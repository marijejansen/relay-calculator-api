<?xml version="1.0" encoding="ISO-8859-1"?>
<LENEX version="2.0">
 <CONSTRUCTOR name="KNZB masters db" version="1.0">
  <CONTACT name="Grove" email="zwemgrove@kpnmail.nl" />
 </CONSTRUCTOR>
 <RECORDLISTS>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="20" agemax="24" />
   <RECORDS>
    <RECORD swimtime="00:00:26.20">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <ATHLETE firstname="Saranda" nameprefix="" lastname="Hofstra" gender="F" nation="NED" CLUB="KSN (SG)" birthdate="1997-03-30" />
    </RECORD>
    <RECORD swimtime="00:00:57.26">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Tamara" nameprefix="" lastname="Grove" gender="F" nation="NED" CLUB="De Dolfijn" birthdate="1996-10-02" />
    </RECORD>
    <RECORD swimtime="00:02:04.07">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Tamara" nameprefix="" lastname="Grove" gender="F" nation="NED" CLUB="De Dolfijn" birthdate="1996-10-02" />
    </RECORD>
    <RECORD swimtime="00:04:20.22">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Madelon" nameprefix="" lastname="Dijkstra" gender="F" nation="NED" CLUB="ZPCH" birthdate="1997-11-04" />
    </RECORD>
    <RECORD swimtime="00:08:53.47">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Madelon" nameprefix="" lastname="Dijkstra" gender="F" nation="NED" CLUB="ZPCH" birthdate="1997-11-04" />
    </RECORD>
    <RECORD swimtime="00:16:49.30">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-23" nation="NED" />
     <ATHLETE firstname="Madelon" nameprefix="" lastname="Dijkstra" gender="F" nation="NED" CLUB="ZPCH" birthdate="1997-11-04" />
    </RECORD>
    <RECORD swimtime="00:00:28.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <ATHLETE firstname="Britta" nameprefix="" lastname="Koehorst" gender="F" nation="NED" CLUB="WVZ" birthdate="2003-05-03" />
    </RECORD>
    <RECORD swimtime="00:01:02.93">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <ATHLETE firstname="Saranda" nameprefix="" lastname="Hofstra" gender="F" nation="NED" CLUB="KSN (SG)" birthdate="1997-03-30" />
    </RECORD>
    <RECORD swimtime="00:02:17.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Almere-Poort" date="2018-11-18" nation="NED" />
     <ATHLETE firstname="Jamilla" nameprefix="van" lastname="Veen" gender="F" nation="NED" CLUB="Zwemvereniging Hoogland" birthdate="1996-07-24" />
    </RECORD>
    <RECORD swimtime="00:00:31.65">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <ATHLETE firstname="Anne Louise" nameprefix="" lastname="Palmans" gender="F" nation="NED" CLUB="WVZ" birthdate="2000-07-27" />
    </RECORD>
    <RECORD swimtime="00:01:10.22">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <ATHLETE firstname="Anne Louise" nameprefix="" lastname="Palmans" gender="F" nation="NED" CLUB="WVZ" birthdate="2000-07-27" />
    </RECORD>
    <RECORD swimtime="00:02:39.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Chantal" nameprefix="van der" lastname="Horst" gender="F" nation="NED" CLUB="De Meer" birthdate="1994-01-08" />
    </RECORD>
    <RECORD swimtime="00:00:27.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <ATHLETE firstname="Britta" nameprefix="" lastname="Koehorst" gender="F" nation="NED" CLUB="WVZ" birthdate="2003-05-03" />
    </RECORD>
    <RECORD swimtime="00:01:03.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Nijverdal" date="2013-01-27" nation="NED" />
     <ATHLETE firstname="Chantal" nameprefix="" lastname="Nap" gender="F" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1989-04-08" />
    </RECORD>
    <RECORD swimtime="00:02:18.46">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2014-01-25" nation="NED" />
     <ATHLETE firstname="Lisa" nameprefix="" lastname="Dreesens" gender="F" nation="NED" CLUB="PSV" birthdate="1991-10-05" />
    </RECORD>
    <RECORD swimtime="00:01:02.33">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <ATHLETE firstname="Britta" nameprefix="" lastname="Koehorst" gender="F" nation="NED" CLUB="WVZ" birthdate="2003-05-03" />
    </RECORD>
    <RECORD swimtime="00:02:20.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <ATHLETE firstname="Anne Louise" nameprefix="" lastname="Palmans" gender="F" nation="NED" CLUB="WVZ" birthdate="2000-07-27" />
    </RECORD>
    <RECORD swimtime="00:04:56.90">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Madelon" nameprefix="" lastname="Dijkstra" gender="F" nation="NED" CLUB="ZPCH" birthdate="1997-11-04" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:25.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-12-23" nation="NED" />
     <ATHLETE firstname="Clarissa" nameprefix="van" lastname="Rheenen" gender="F" nation="NED" CLUB="PSV" birthdate="1991-06-26" />
    </RECORD>
    <RECORD swimtime="00:00:54.92">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Marjolein" nameprefix="" lastname="Delno" gender="F" nation="NED" CLUB="VZC" birthdate="1994-03-17" />
    </RECORD>
    <RECORD swimtime="00:01:57.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" CLUB="De Dolfijn" birthdate="1998-01-29" />
    </RECORD>
    <RECORD swimtime="00:04:13.71">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" CLUB="De Dolfijn" birthdate="1998-01-29" />
    </RECORD>
    <RECORD swimtime="00:09:17.98">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vlissingen" date="2005-03-06" nation="NED" />
     <ATHLETE firstname="Maartje" nameprefix="van" lastname="Keulen" gender="F" nation="NED" CLUB="SBC2000" birthdate="1980-01-01" />
    </RECORD>
    <RECORD swimtime="00:17:53.76">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Winterswijk" date="2005-01-23" nation="NED" />
     <ATHLETE firstname="Elvira" nameprefix="" lastname="Jonkers" gender="F" nation="NED" CLUB="TriVia" birthdate="1979-10-31" />
    </RECORD>
    <RECORD swimtime="00:00:30.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Dronten" date="2017-06-03" nation="NED" />
     <ATHLETE firstname="Elinore" nameprefix="de" lastname="Jong" gender="F" nation="NED" CLUB="The Hague Swimming (SG)" birthdate="1989-04-23" />
    </RECORD>
    <RECORD swimtime="00:01:03.84">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" CLUB="De Dolfijn" birthdate="1998-01-29" />
    </RECORD>
    <RECORD swimtime="00:02:10.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" CLUB="De Dolfijn" birthdate="1998-01-29" />
    </RECORD>
    <RECORD swimtime="00:00:32.37">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2018-12-02" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Brouwer" gender="F" nation="NED" CLUB="SwimGym" birthdate="1991-03-02" />
    </RECORD>
    <RECORD swimtime="00:01:12.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Yvon" nameprefix="" lastname="Versteeg" gender="F" nation="NED" CLUB="De Veene" birthdate="1992-03-31" />
    </RECORD>
    <RECORD swimtime="00:02:37.59">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Yvon" nameprefix="" lastname="Versteeg" gender="F" nation="NED" CLUB="De Veene" birthdate="1992-03-31" />
    </RECORD>
    <RECORD swimtime="00:00:26.14">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Elinore" nameprefix="de" lastname="Jong" gender="F" nation="NED" CLUB="The Hague Swimming (SG)" birthdate="1989-04-23" />
    </RECORD>
    <RECORD swimtime="00:01:00.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Dronten" date="2017-06-03" nation="NED" />
     <ATHLETE firstname="Elinore" nameprefix="de" lastname="Jong" gender="F" nation="NED" CLUB="The Hague Swimming (SG)" birthdate="1989-04-23" />
    </RECORD>
    <RECORD swimtime="00:02:19.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Vlissingen" date="2005-03-06" nation="NED" />
     <ATHLETE firstname="Sandra" nameprefix="" lastname="Temmerman" gender="F" nation="NED" CLUB="SBC2000" birthdate="1980-01-09" />
    </RECORD>
    <RECORD swimtime="00:01:04.71">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Yvon" nameprefix="" lastname="Versteeg" gender="F" nation="NED" CLUB="De Veene" birthdate="1992-03-31" />
    </RECORD>
    <RECORD swimtime="00:02:21.39">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Inge" nameprefix="" lastname="Arts" gender="F" nation="NED" CLUB="Merlet" birthdate="1992-05-29" />
    </RECORD>
    <RECORD swimtime="00:05:05.12">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <ATHLETE firstname="Inge" nameprefix="" lastname="Arts" gender="F" nation="NED" CLUB="Merlet" birthdate="1992-05-29" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:24.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Derby" date="2023-11-26" nation="GBR" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Hopkin" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:52.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Derby" date="2023-11-25" nation="GBR" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Hopkin" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:57.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:04:13.71">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:08:57.67">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gau Algesheim" date="2009-01-17" nation="GER" />
     <ATHLETE firstname="Susanne" nameprefix="" lastname="Keller" gender="F" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:16:47.66">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gau Algesheim" date="2009-01-17" nation="GER" />
     <ATHLETE firstname="Susanne" nameprefix="" lastname="Keller" gender="F" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:00:28.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2023-10-29" nation="GBR" />
     <ATHLETE firstname="Georgina" nameprefix="" lastname="Pryor" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:01.23">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Poznan" date="2022-12-17" nation="POL" />
     <ATHLETE firstname="Gabriela" nameprefix="" lastname="Wojtowicz" gender="F" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:02:10.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:30.50">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Ceska Lipa" date="2014-06-08" nation="CZE" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Chocova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:06.83">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Ceska Lipa" date="2014-06-07" nation="CZE" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Chocova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:30.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2009-10-24" nation="GBR" />
     <ATHLETE firstname="Katie" nameprefix="" lastname="Henderson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:26.14">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Elinore" nameprefix="de" lastname="Jong" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:58.98">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="2023-10-29" nation="GBR" />
     <ATHLETE firstname="Georgina" nameprefix="" lastname="Pryor" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:17.11">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Hamburg" date="2017-11-11" nation="GER" />
     <ATHLETE firstname="Lisa" nameprefix="" lastname="Stamm" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:02.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Ceska Lipa" date="2014-06-08" nation="CZE" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Chocova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:17.54">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Palma de Mallorca" date="2014-02-21" nation="ESP" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Markova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:04:44.98">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Recklinghausen" date="2015-09-27" nation="GER" />
     <ATHLETE firstname="Katarzyna" nameprefix="" lastname="Baranowska" gender="F" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:24.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-10-27" nation="" />
     <ATHLETE firstname="Rebecca" nameprefix="" lastname="Guy" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:54.44">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-11-16" nation="" />
     <ATHLETE firstname="Yayoi" nameprefix="" lastname="Matsumoto" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:57.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:04:13.71">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:08:51.18">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="1996-03-31" nation="" />
     <ATHLETE firstname="Sheila" nameprefix="" lastname="Taormina" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:16:36.07">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="1996-03-31" nation="" />
     <ATHLETE firstname="Sheila" nameprefix="" lastname="Taormina" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:27.88">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2015-06-14" nation="" />
     <ATHLETE firstname="Yurie" nameprefix="" lastname="Oga" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:00.63">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2015-10-05" nation="" />
     <ATHLETE firstname="Yurie" nameprefix="" lastname="Oga" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:10.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:30.50">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Ceska Lipa" date="2014-06-08" nation="CZE" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Chocova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:06.83">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Ceska Lipa" date="2014-06-07" nation="CZE" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Chocova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:28.33">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-03-21" nation="" />
     <ATHLETE firstname="Satori" nameprefix="" lastname="Hosokoshi" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:26.14">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Elinore" nameprefix="de" lastname="Jong" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:58.11">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2015-12-12" nation="" />
     <ATHLETE firstname="Claire" nameprefix="" lastname="Donahue" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:09.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2010-05-08" nation="" />
     <ATHLETE firstname="Yuko" nameprefix="" lastname="Nakanishi" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:01.79">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-01-26" nation="" />
     <ATHLETE firstname="Masako" nameprefix="" lastname="Kuroki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:17.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2006-04-23" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:04:44.98">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-09-27" nation="" />
     <ATHLETE firstname="Katarzyna" nameprefix="" lastname="Baranowska" gender="F" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:26.41">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Saskia" nameprefix="de" lastname="Klerk" gender="F" nation="NED" CLUB="GoSwim" birthdate="1990-11-29" />
    </RECORD>
    <RECORD swimtime="00:00:57.02">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <ATHLETE firstname="Pauline" nameprefix="" lastname="Gouwens" gender="F" nation="NED" CLUB="DWK" birthdate="1984-11-23" />
    </RECORD>
    <RECORD swimtime="00:02:05.69">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" CLUB="WVZ" birthdate="1993-11-05" />
    </RECORD>
    <RECORD swimtime="00:04:28.31">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" CLUB="WVZ" birthdate="1993-11-05" />
    </RECORD>
    <RECORD swimtime="00:09:16.42">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" CLUB="WVZ" birthdate="1993-11-05" />
    </RECORD>
    <RECORD swimtime="00:18:06.33">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Emmeloord" date="2006-01-22" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Het Y" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:00:30.94">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Evy" nameprefix="" lastname="Witlox" gender="F" nation="NED" CLUB="DWT" birthdate="1988-08-28" />
    </RECORD>
    <RECORD swimtime="00:01:06.30">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <ATHLETE firstname="Evy" nameprefix="" lastname="Witlox" gender="F" nation="NED" CLUB="DWT" birthdate="1988-08-28" />
    </RECORD>
    <RECORD swimtime="00:02:20.26">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" CLUB="WVZ" birthdate="1993-11-05" />
    </RECORD>
    <RECORD swimtime="00:00:33.03">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2015-01-24" nation="NED" />
     <ATHLETE firstname="Karin" nameprefix="" lastname="Hidding" gender="F" nation="NED" CLUB="De Dinkel" birthdate="1984-01-08" />
    </RECORD>
    <RECORD swimtime="00:01:12.74">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1988-07-28" />
    </RECORD>
    <RECORD swimtime="00:02:41.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1988-07-28" />
    </RECORD>
    <RECORD swimtime="00:00:27.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2015-01-23" nation="NED" />
     <ATHLETE firstname="Pauline" nameprefix="" lastname="Gouwens" gender="F" nation="NED" CLUB="DWK" birthdate="1984-11-23" />
    </RECORD>
    <RECORD swimtime="00:01:03.12">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2014-01-24" nation="NED" />
     <ATHLETE firstname="Pauline" nameprefix="" lastname="Gouwens" gender="F" nation="NED" CLUB="DWK" birthdate="1984-11-23" />
    </RECORD>
    <RECORD swimtime="00:02:24.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Winterswijk" date="2002-05-04" nation="NED" />
     <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" CLUB="AZ&amp;PC" birthdate="1970-07-01" />
    </RECORD>
    <RECORD swimtime="00:01:07.72">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Winterswijk" date="2002-05-03" nation="NED" />
     <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" CLUB="AZ&amp;PC" birthdate="1970-07-01" />
    </RECORD>
    <RECORD swimtime="00:02:26.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Winterswijk" date="2002-05-05" nation="NED" />
     <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" CLUB="AZ&amp;PC" birthdate="1970-07-01" />
    </RECORD>
    <RECORD swimtime="00:05:03.27">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Marlijn" nameprefix="" lastname="Hendriksen" gender="F" nation="NED" CLUB="Hieronymus" birthdate="1988-08-16" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:24.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-28" nation="GBR" />
     <ATHLETE firstname="Rebecca" nameprefix="" lastname="Guy" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:55.11">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Bordeaux" date="2009-01-25" nation="FRA" />
     <ATHLETE firstname="Alena" nameprefix="" lastname="Popchanka" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:02.03">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2017-10-27" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:04:14.56">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2017-10-28" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:42.57">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2017-10-29" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:17:02.39">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2018-10-26" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:28.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Esbjerg" date="2006-03-25" nation="DEN" />
     <ATHLETE firstname="Mette" nameprefix="" lastname="Jacobsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:01:02.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Esbjerg" date="2006-03-26" nation="DEN" />
     <ATHLETE firstname="Mette" nameprefix="" lastname="Jacobsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:02:13.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2017-10-28" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:31.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Ceska Lipa" date="2016-11-13" nation="CZE" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Chocova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:08.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Ceska Lipa" date="2016-11-12" nation="CZE" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Chocova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:32.71">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2018-10-27" nation="GBR" />
     <ATHLETE firstname="Georgina" nameprefix="" lastname="Heyn" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:26.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="2023-10-27" nation="GBR" />
     <ATHLETE firstname="Rebecca" nameprefix="" lastname="Guy" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:59.82">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Kazan" date="2016-11-20" nation="RUS" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Polyakova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:19.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Lecco" date="2004-03-27" nation="ITA" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Bianzani" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:03.31">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Ceska Lipa" date="2016-11-13" nation="CZE" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Chocova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:16.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Epinal" date="2016-01-31" nation="FRA" />
     <ATHLETE firstname="Sophie" nameprefix="de" lastname="Ronchi" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:50.66">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="St. Petersburg" date="2014-11-28" nation="RUS" />
     <ATHLETE firstname="Natalia" nameprefix="" lastname="Vinokourenkova" gender="F" nation="RUS" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:25.17">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-11-29" nation="" />
     <ATHLETE firstname="Svetlana" nameprefix="" lastname="Kniaginina" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:54.75">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2012-10-13" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Erndl" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:00.73">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-11-14" nation="" />
     <ATHLETE firstname="Veronica" nameprefix="" lastname="Balsano" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:04:14.56">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-10-28" nation="" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:38.58">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-12-04" nation="" />
     <ATHLETE firstname="Dawn" nameprefix="" lastname="Heckman" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:16:26.93">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-12-02" nation="" />
     <ATHLETE firstname="Dawn" nameprefix="" lastname="Heckman" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:27.43">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2009-04-19" nation="" />
     <ATHLETE firstname="Mai" nameprefix="" lastname="Nakamura" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:00.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2010-03-07" nation="" />
     <ATHLETE firstname="Kana" nameprefix="" lastname="Yamaguchi" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:11.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2012-04-21" nation="" />
     <ATHLETE firstname="Kana" nameprefix="" lastname="Yamaguchi" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:31.35">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2015-11-29" nation="" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:06.98">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-04-17" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:26.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2009-04-18" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:26.67">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-03-18" nation="" />
     <ATHLETE firstname="Masako" nameprefix="" lastname="Ida" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:59.82">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Kazan" date="2016-11-20" nation="RUS" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Polyakova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:13.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2008-05-25" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:02.52">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2012-10-13" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Erndl" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:13.41">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-11-14" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:04:45.07">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2010-04-17" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:27.27">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Anneloes" nameprefix="" lastname="Peulen" gender="F" nation="NED" CLUB="Nuenen" birthdate="1985-04-25" />
    </RECORD>
    <RECORD swimtime="00:00:59.65">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Pauline" nameprefix="" lastname="Gouwens" gender="F" nation="NED" CLUB="DWK" birthdate="1984-11-23" />
    </RECORD>
    <RECORD swimtime="00:02:11.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:04:37.34">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Grootebroek" date="2017-05-21" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:09:34.16">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Winterswijk" date="2008-04-02" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Het Y" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:18:16.12">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Winterswijk" date="2008-05-04" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Het Y" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:00:31.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1985-09-29" />
    </RECORD>
    <RECORD swimtime="00:01:09.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Maastricht" date="2017-01-20" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:32.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Schouten" gender="F" nation="NED" CLUB="MZ&amp;PC" birthdate="1987-09-08" />
    </RECORD>
    <RECORD swimtime="00:00:34.16">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <ATHLETE firstname="Loes" nameprefix="" lastname="Zanderink" gender="F" nation="NED" CLUB="SwimGym" birthdate="1988-11-23" />
    </RECORD>
    <RECORD swimtime="00:01:14.67">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2023-11-26" nation="NED" />
     <ATHLETE firstname="Loes" nameprefix="" lastname="Zanderink" gender="F" nation="NED" CLUB="SwimGym" birthdate="1988-11-23" />
    </RECORD>
    <RECORD swimtime="00:02:49.21">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="DAW" birthdate="1982-04-05" />
    </RECORD>
    <RECORD swimtime="00:00:28.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <ATHLETE firstname="Pauline" nameprefix="" lastname="Gouwens" gender="F" nation="NED" CLUB="DWK" birthdate="1984-11-23" />
    </RECORD>
    <RECORD swimtime="00:01:06.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:30.69">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Maastricht" date="2017-01-20" nation="NED" />
     <ATHLETE firstname="Roos" nameprefix="van" lastname="Esch" gender="F" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1982-07-17" />
    </RECORD>
    <RECORD swimtime="00:01:08.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:29.83">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Maastricht" date="2017-01-20" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:05:28.27">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <ATHLETE firstname="Roos" nameprefix="van" lastname="Esch" gender="F" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1982-07-17" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:25.91">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sori" date="2015-01-18" nation="ITA" />
     <ATHLETE firstname="Olessia" nameprefix="" lastname="Bourova" gender="F" nation="ita" />
    </RECORD>
    <RECORD swimtime="00:00:57.12">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2010-10-29" nation="GBR" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Roca" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:04.92">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Pontevedra" date="2015-02-20" nation="ESP" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Roca" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:04:19.96">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Stockport" date="2023-07-15" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:50.76">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Carlisle" date="2020-01-31" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:17:26.96">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Blackpool" date="2018-02-24" nation="GBR" />
     <ATHLETE firstname="Emma" nameprefix="" lastname="Wills" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:29.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Norwich" date="2009-05-16" nation="GBR" />
     <ATHLETE firstname="Zoe" nameprefix="" lastname="Cray" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:03.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2009-10-24" nation="GBR" />
     <ATHLETE firstname="Zoe" nameprefix="" lastname="Cray" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:17.11">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2023-10-29" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:30.96">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Funchal" date="2023-11-20" nation="POR" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Weber" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:08.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Ceska Lipa" date="2023-11-11" nation="CZE" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Weber" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:35.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Twist" date="2017-05-21" nation="GER" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:27.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Funchal" date="2023-11-23" nation="POR" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Weber" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:02.92">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Saransk" date="2021-11-13" nation="RUS" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Polyakova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:20.92">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Vikt�ria" nameprefix="" lastname="H�den-Felf�ldi" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:01:02.76">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Funchal" date="2023-11-19" nation="POR" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Weber" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:20.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2018-11-17" nation="RUS" />
     <ATHLETE firstname="Natalia" nameprefix="" lastname="Vinokourenkova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:05:00.31">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2018-11-16" nation="RUS" />
     <ATHLETE firstname="Natalia" nameprefix="" lastname="Vinokourenkova" gender="F" nation="RUS" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:25.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2006-12-03" nation="" />
     <ATHLETE firstname="Dara" nameprefix="" lastname="Torres" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:54.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2006-12-03" nation="" />
     <ATHLETE firstname="Dara" nameprefix="" lastname="Torres" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:03.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2012-03-25" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:04:19.96">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-07-15" nation="" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:50.76">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2020-01-31" nation="" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:16:52.94">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-09-27" nation="" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:27.63">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2016-11-13" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:00.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-11-19" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:13.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2013-11-16" nation="" />
     <ATHLETE firstname="Kana" nameprefix="" lastname="Ohashi" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:31.25">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-10-08" nation="USA" />
     <ATHLETE firstname="Danielle" nameprefix="" lastname="Herrmann" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:08.59">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-10-08" nation="USA" />
     <ATHLETE firstname="Danielle" nameprefix="" lastname="Herrmann" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:30.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2012-03-10" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:27.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-10-08" nation="USA" />
     <ATHLETE firstname="Danielle" nameprefix="" lastname="Herrmann" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:01.31">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-07-25" nation="BRA" />
     <ATHLETE firstname="Carolina" nameprefix="" lastname="Athayde" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:02:14.46">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-07-24" nation="" />
     <ATHLETE firstname="Carolina" nameprefix="" lastname="Athayde" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:01:03.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2012-03-10" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:17.69">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2012-11-18" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:04:52.85">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="1997-12-14" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:27.72">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:01:00.19">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:11.83">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwijndrecht" date="2023-12-16" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:04:42.74">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-25" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:09:33.98">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-24" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:18:11.24">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-26" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:00:32.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwolle" date="2014-01-25" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:01:09.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Breda" date="2015-11-08" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:02:32.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Nijlen" date="2016-03-19" nation="BEL" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:00:35.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Oss" date="2022-09-25" nation="NED" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="DAW" birthdate="1982-04-05" />
    </RECORD>
    <RECORD swimtime="00:01:18.24">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:49.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="DAW" birthdate="1982-04-05" />
    </RECORD>
    <RECORD swimtime="00:00:29.40">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:01:06.94">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Papendrecht" date="2022-10-09" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:33.44">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Vlaardingen" date="2010-01-22" nation="NED" />
     <ATHLETE firstname="Anita" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="DIO" birthdate="1969-10-12" />
    </RECORD>
    <RECORD swimtime="00:01:07.94">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:31.71">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Oss" date="2022-09-25" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:05:30.28">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2015-01-24" nation="NED" />
     <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" CLUB="PSV" birthdate="1975-03-04" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:26.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Essen" date="2021-11-27" nation="GER" />
     <ATHLETE firstname="Katja" nameprefix="" lastname="Otto" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:58.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Lappeenrannan" date="2017-03-18" nation="FIN" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:02:07.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Jersey" date="2014-09-13" nation="GBR" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:04:24.42">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Jersey" date="2014-09-13" nation="GBR" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:08:55.34">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-24" nation="NED" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:17:01.66">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Wigan" date="2015-02-22" nation="GBR" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:29.84">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Newmarket" date="2014-10-04" nation="GBR" />
     <ATHLETE firstname="Zoe" nameprefix="" lastname="Cray" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:03.22">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Salo" date="2018-03-24" nation="FIN" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:02:21.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2012-10-26" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:31.81">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rostock" date="2022-11-20" nation="GER" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:10.16">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Baunatal" date="2022-11-05" nation="GER" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:32.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Baunatal" date="2022-11-05" nation="GER" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:28.33">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2015-02-14" nation="ITA" />
     <ATHLETE firstname="Roberta" nameprefix="" lastname="Crescentini" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:03.76">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Kastrup" date="2015-11-07" nation="DEN" />
     <ATHLETE firstname="Sophia" nameprefix="" lastname="Skou" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:02:24.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Malm�" date="2018-10-12" nation="SWE" />
     <ATHLETE firstname="Sophia" nameprefix="" lastname="Skou" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:01:04.32">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Espoo" date="2018-01-13" nation="FIN" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:02:24.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Mansea" date="2021-04-17" nation="ESP" />
     <ATHLETE firstname="Mirea" nameprefix="" lastname="Garcia" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:05:06.66">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Mansea" date="2021-04-17" nation="ESP" />
     <ATHLETE firstname="Mirea" nameprefix="" lastname="Garcia" gender="F" nation="ESP" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:26.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-12-14" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:57.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-12-14" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:05.26">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2003-12-14" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:21.75">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2003-12-14" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:08:55.34">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-24" nation="NED" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:16:50.92">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-12-01" nation="" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-01-14" nation="" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:01:03.22">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-03-24" nation="" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:02:17.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-05-27" nation="" />
     <ATHLETE firstname="Kana" nameprefix="" lastname="Morihisa" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:32.16">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-12-02" nation="" />
     <ATHLETE firstname="Katie" nameprefix="" lastname="Glenn" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:09.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2015-12-05" nation="" />
     <ATHLETE firstname="Cynthia" nameprefix="" lastname="Lewis" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:32.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2008-11-16" nation="" />
     <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2013-03-16" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:01.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2009-11-21" nation="" />
     <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:20.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2006-11-19" nation="" />
     <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:04.19">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-10-10" nation="" />
     <ATHLETE firstname="Lisa" nameprefix="" lastname="Blackburn" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:19.21">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2007-12-02" nation="" />
     <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:00.82">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2002-11-24" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:27.91">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2015-01-25" nation="NED" />
     <ATHLETE firstname="Monique" nameprefix="" lastname="Tuijp" gender="F" nation="NED" CLUB="WZ&amp;PC Purmerend" birthdate="1969-01-28" />
    </RECORD>
    <RECORD swimtime="00:01:02.16">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Lelystad" date="2014-12-20" nation="NED" />
     <ATHLETE firstname="Monique" nameprefix="" lastname="Tuijp" gender="F" nation="NED" CLUB="WZ&amp;PC Purmerend" birthdate="1969-01-28" />
    </RECORD>
    <RECORD swimtime="00:02:07.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" CLUB="PSV" birthdate="1973-11-06" />
    </RECORD>
    <RECORD swimtime="00:04:47.60">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Leiden" date="2024-01-21" nation="NED" />
     <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" CLUB="PSV" birthdate="1975-03-04" />
    </RECORD>
    <RECORD swimtime="00:09:49.67">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="De Otters Het Gooi" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:18:48.97">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-23" nation="NED" />
     <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" CLUB="PSV" birthdate="1975-03-04" />
    </RECORD>
    <RECORD swimtime="00:00:33.38">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Edith" nameprefix="" lastname="Janssen-Koolen" gender="F" nation="NED" CLUB="TRB-RES" birthdate="1973-01-10" />
    </RECORD>
    <RECORD swimtime="00:01:10.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:02:32.98">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1972-03-08" />
    </RECORD>
    <RECORD swimtime="00:00:34.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Maastricht" date="2017-01-20" nation="NED" />
     <ATHLETE firstname="Marjo" nameprefix="" lastname="Goelema-Koek" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1969-01-02" />
    </RECORD>
    <RECORD swimtime="00:01:18.62">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <ATHLETE firstname="Marjo" nameprefix="" lastname="Goelema-Koek" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1969-01-02" />
    </RECORD>
    <RECORD swimtime="00:02:54.04">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2014-01-25" nation="NED" />
     <ATHLETE firstname="Annette" nameprefix="" lastname="Wijnja-Visser" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1967-01-30" />
    </RECORD>
    <RECORD swimtime="00:00:30.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Papendrecht" date="2016-01-24" nation="NED" />
     <ATHLETE firstname="Ingrid" nameprefix="" lastname="Boot-de Groot" gender="F" nation="NED" CLUB="De Aalscholver" birthdate="1970-08-08" />
    </RECORD>
    <RECORD swimtime="00:01:10.01">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Jeanne" nameprefix="" lastname="Petit" gender="F" nation="NED" CLUB="De Dinkel" birthdate="1970-02-13" />
    </RECORD>
    <RECORD swimtime="00:02:38.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2020-01-04" nation="NED" />
     <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" CLUB="PSV" birthdate="1975-03-04" />
    </RECORD>
    <RECORD swimtime="00:01:11.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:02:35.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Emmeloord" date="2019-03-16" nation="NED" />
     <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1972-03-08" />
    </RECORD>
    <RECORD swimtime="00:05:32.35">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Leiden" date="2020-02-23" nation="NED" />
     <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" CLUB="PSV" birthdate="1975-03-04" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:26.37">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Paris" date="2013-05-18" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:58.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Paris" date="2014-03-29" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:07.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:04:37.53">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Trondheim" date="2016-04-09" nation="NOR" />
     <ATHLETE firstname="Merete" nameprefix="" lastname="L�vberg" gender="F" nation="NOR" />
    </RECORD>
    <RECORD swimtime="00:09:25.12">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Copenhagen" date="2010-01-16" nation="DEN" />
     <ATHLETE firstname="Susanna" nameprefix="" lastname="Ros�n" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:17:57.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Lodi" date="2016-02-13" nation="ITA" />
     <ATHLETE firstname="Valeria" nameprefix="" lastname="Vergani" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:29.52">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Espoo" date="2020-01-11" nation="FIN" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:01:05.76">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2018-10-26" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:20.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2016-10-28" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:33.56">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2009-01-11" nation="ITA" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:11.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Desenzano" date="2009-01-25" nation="ITA" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:37.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Desenzano" date="2009-01-25" nation="ITA" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:28.79">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2020-02-16" nation="ITA" />
     <ATHLETE firstname="Roberta" nameprefix="" lastname="Crescentini" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:05.83">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2016-04-03" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Soro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:26.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Flensburg" date="2014-02-15" nation="GER" />
     <ATHLETE firstname="Barbara" nameprefix="" lastname="Kehbein" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:06.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="S�dert�lje" date="2013-03-16" nation="SWE" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Hammar" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:02:26.98">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Vienna" date="2022-04-02" nation="AUT" />
     <ATHLETE firstname="Smiljana" nameprefix="" lastname="Marinovic" gender="F" nation="CRO" />
    </RECORD>
    <RECORD swimtime="00:05:17.83">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Espoo" date="2018-04-20" nation="FIN" />
     <ATHLETE firstname="Satu" nameprefix="" lastname="Rahkonen" gender="F" nation="FIN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:26.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-10-13" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:57.89">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-09-12" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:05.94">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2007-12-02" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:24.86">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-08-01" nation="" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:01.09">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-01-28" nation="USA" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:01.27">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-01-28" nation="USA" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:29.52">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2020-01-11" nation="" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:01:04.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2009-02-27" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:18.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2009-02-26" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:33.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-07-16" nation="" />
     <ATHLETE firstname="Linley" nameprefix="" lastname="Frame" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:10.63">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-07-16" nation="" />
     <ATHLETE firstname="Linley" nameprefix="" lastname="Frame" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:02:34.77">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-12-02" nation="" />
     <ATHLETE firstname="Gabrielle" nameprefix="" lastname="Rose" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.53">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-10-15" nation="" />
     <ATHLETE firstname="Yuriko" nameprefix="" lastname="Ikeda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:03.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2010-11-20" nation="" />
     <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:23.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2009-12-13" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:05.61">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-02-26" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:19.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-12-02" nation="" />
     <ATHLETE firstname="Gabrielle" nameprefix="" lastname="Rose" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:00.29">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-02-27" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:28.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Monique" nameprefix="" lastname="Tuijp" gender="F" nation="NED" CLUB="WZ&amp;PC Purmerend" birthdate="1969-01-28" />
    </RECORD>
    <RECORD swimtime="00:01:02.83">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:02:17.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:04:40.53">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:09:38.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2022-09-24" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:18:14.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2022-09-24" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:00:33.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Maastricht" date="2022-12-29" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:01:11.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kapelle" date="2022-04-03" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:02:41.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwolle" date="2014-01-26" nation="NED" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Cromjongh" gender="F" nation="NED" CLUB="De Zwoer" birthdate="1964-03-17" />
    </RECORD>
    <RECORD swimtime="00:00:35.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Marjo" nameprefix="" lastname="Goelema-Koek" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1969-01-02" />
    </RECORD>
    <RECORD swimtime="00:01:19.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" CLUB="PSV" birthdate="1970-03-02" />
    </RECORD>
    <RECORD swimtime="00:02:55.02">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" CLUB="PSV" birthdate="1970-03-02" />
    </RECORD>
    <RECORD swimtime="00:00:31.25">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Jeanne" nameprefix="" lastname="Petit" gender="F" nation="NED" CLUB="PSV" birthdate="1970-02-13" />
    </RECORD>
    <RECORD swimtime="00:01:09.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Oss" date="2022-09-25" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:02:39.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Vlissingen" date="2009-01-23" nation="NED" />
     <ATHLETE firstname="Mathilde" nameprefix="" lastname="Vink" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1958-12-12" />
    </RECORD>
    <RECORD swimtime="00:01:12.64">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Oss" date="2022-09-25" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:02:34.81">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Oss" date="2022-09-25" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:05:45.52">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Almere-Poort" date="2023-03-12" nation="NED" />
     <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1970-07-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:26.27">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rennes" date="2015-03-27" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:58.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Montlugon" date="2015-01-25" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:11.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Dunkerque" date="2017-03-23" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:39.14">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Torino" date="2023-12-08" nation="ITA" />
     <ATHLETE firstname="Tiziana" nameprefix="" lastname="Papandrea" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:09:38.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2022-09-24" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:18:14.50">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2022-09-24" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:31.16">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rennes" date="2015-03-28" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:06.52">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2022-10-28" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:26.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2022-10-30" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:34.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Trento" date="2012-03-18" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Soro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:13.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="London" date="2022-07-10" nation="GBR" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:41.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:29.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="J�nk�ping" date="2018-03-25" nation="SWE" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Hammar" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:01:06.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Brescia" date="2016-04-03" nation="ITA" />
     <ATHLETE firstname="Daniela" nameprefix="de" lastname="Ponti" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:28.69">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Riccione" date="2018-02-25" nation="ITA" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:07.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Kastrup" date="2015-11-07" nation="DEN" />
     <ATHLETE firstname="Anette" nameprefix="" lastname="Philipsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:02:30.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Derby" date="2023-11-25" nation="GBR" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:05:23.74">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Stockport" date="2023-07-15" nation="GBR" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:26.27">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-03-27" nation="" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:58.12">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-10-15" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:10.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-12-06" nation="" />
     <ATHLETE firstname="Suzanne" nameprefix="" lastname="Heim-Bowen" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:33.86">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-17" nation="" />
     <ATHLETE firstname="Alison" nameprefix="" lastname="Zamanian" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:23.30">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-16" nation="" />
     <ATHLETE firstname="Alison" nameprefix="" lastname="Zamanian" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:47.04">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-01-29" nation="" />
     <ATHLETE firstname="Alison" nameprefix="" lastname="Zamanian" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:30.27">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2015-12-13" nation="" />
     <ATHLETE firstname="Leslie" nameprefix="" lastname="Livingston" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:05.89">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2014-03-08" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:22.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2014-03-08" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:33.96">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2012-11-24" nation="" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:13.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-07-10" nation="" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:41.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-10-29" nation="" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:28.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-06-17" nation="" />
     <ATHLETE firstname="Susan" nameprefix="" lastname="O'Neill" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:06.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-09-25" nation="" />
     <ATHLETE firstname="Yuriko" nameprefix="" lastname="Ikeda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:28.08">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2011-05-08" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:07.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-10-15" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:27.39">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-11-17" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:10.96">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2014-09-26" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:29.31">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Steenwijk" date="2022-04-02" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:01:05.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwijndrecht" date="2022-04-09" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:02:27.48">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC Woerden" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:05:13.76">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gorinchem" date="2018-03-03" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC Woerden" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:11:00.20">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <ATHLETE firstname="Wilna" nameprefix="" lastname="Heijman-Hartkamp" gender="F" nation="NED" CLUB="Steenwijk 1934" birthdate="1964-05-03" />
    </RECORD>
    <RECORD swimtime="00:21:02.61">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-19" nation="NED" />
     <ATHLETE firstname="Irene" nameprefix="van der" lastname="Laan" gender="F" nation="NED" CLUB="ZV De Bron" birthdate="1960-12-27" />
    </RECORD>
    <RECORD swimtime="00:00:35.33">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Steenwijk" date="2022-04-02" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:01:16.63">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwijndrecht" date="2022-04-09" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:02:42.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Cromjongh" gender="F" nation="NED" CLUB="De Zwoer" birthdate="1964-03-17" />
    </RECORD>
    <RECORD swimtime="00:00:38.31">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2024-01-06" nation="NED" />
     <ATHLETE firstname="Jacqueline" nameprefix="" lastname="Tuin" gender="F" nation="NED" CLUB="DAW" birthdate="1966-04-21" />
    </RECORD>
    <RECORD swimtime="00:01:25.19">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwijndrecht" date="2022-04-09" nation="NED" />
     <ATHLETE firstname="Annette" nameprefix="" lastname="Wijnja-Visser" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1967-01-30" />
    </RECORD>
    <RECORD swimtime="00:03:04.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kapelle" date="2022-04-03" nation="NED" />
     <ATHLETE firstname="Annette" nameprefix="" lastname="Wijnja-Visser" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1967-01-30" />
    </RECORD>
    <RECORD swimtime="00:00:31.88">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Steenwijk" date="2022-04-02" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:01:16.67">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Apeldoorn" date="2014-05-18" nation="NED" />
     <ATHLETE firstname="Mathilde" nameprefix="" lastname="Vink" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1958-12-12" />
    </RECORD>
    <RECORD swimtime="00:02:54.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Nijverdal" date="2013-01-26" nation="NED" />
     <ATHLETE firstname="Mathilde" nameprefix="" lastname="Vink" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1958-12-12" />
    </RECORD>
    <RECORD swimtime="00:01:15.58">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC Woerden" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:02:44.47">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Alphen" date="2018-09-15" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC Woerden" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:05:54.23">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2018-02-17" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC Woerden" birthdate="1963-05-15" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:27.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2022-03-11" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:01.71">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2022-03-11" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:17.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Livorno" date="2023-02-26" nation="ITA" />
     <ATHLETE firstname="Daniela" nameprefix="" lastname="Sabatini" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:04:46.77">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Livorno" date="2023-02-25" nation="ITA" />
     <ATHLETE firstname="Daniela" nameprefix="" lastname="Sabatini" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:09:56.06">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Genova" date="2023-02-19" nation="ITA" />
     <ATHLETE firstname="Daniela" nameprefix="" lastname="Sabatini" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:18:53.01">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Lodi" date="2023-02-18" nation="ITA" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Hoag" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:32.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Forli" date="2023-03-12" nation="ITA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:32.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Forli" date="2023-03-12" nation="ITA" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:10.09">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kastrup" date="2022-11-05" nation="DEN" />
     <ATHLETE firstname="Lise" nameprefix="" lastname="Lothe" gender="F" nation="NOR" />
    </RECORD>
    <RECORD swimtime="00:02:32.08">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Riccione" date="2021-11-21" nation="ITA" />
     <ATHLETE firstname="Silvia" nameprefix="" lastname="Parocchi" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:35.15">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Spresiano" date="2017-04-09" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:17.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Viterbo" date="2019-01-26" nation="ITA" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:46.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Viterbo" date="2019-01-27" nation="ITA" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:30.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Milano" date="2023-12-16" nation="ITA" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:08.11">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Milano" date="2023-12-17" nation="ITA" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:32.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2023-04-22" nation="ITA" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:12.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Genova" date="2020-02-23" nation="ITA" />
     <ATHLETE firstname="Daniela" nameprefix="de" lastname="Ponti" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:36.92">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Freiburg" date="2019-11-29" nation="GER" />
     <ATHLETE firstname="Susanne" nameprefix="" lastname="Reibel-Oberle" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:05:26.95">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Milano" date="2023-12-17" nation="ITA" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:27.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-03-10" nation="" />
     <ATHLETE firstname="Marie-Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:00.61">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-20" nation="NED" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:13.58">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-02-28" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:04:37.35">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-01-23" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:09:32.63">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-04-23" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:18:01.79">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-04-23" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:00:30.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2016-03-05" nation="" />
     <ATHLETE firstname="Leslie" nameprefix="" lastname="Livingston" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:07.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-07-12" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:25.27">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-08-12" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:35.15">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-04-09" nation="" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:17.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-01-26" nation="" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:46.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-01-27" nation="" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:29.39">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2016-03-05" nation="" />
     <ATHLETE firstname="Leslie" nameprefix="" lastname="Livingston" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:08.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:31.13">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2008-09-14" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:09.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:27.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-01-24" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:15.72">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-11-24" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:30.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-24" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:01:07.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:02:28.92">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Almere-Poort" date="2017-11-19" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:05:22.92">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:11:08.25">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" CLUB="PSV" birthdate="1959-05-28" />
    </RECORD>
    <RECORD swimtime="00:21:25.35">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-23" nation="NED" />
     <ATHLETE firstname="Irene" nameprefix="van der" lastname="Laan" gender="F" nation="NED" CLUB="ZVVS" birthdate="1960-12-27" />
    </RECORD>
    <RECORD swimtime="00:00:37.62">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Nijmegen" date="2016-09-17" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:01:21.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:02:57.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:00:41.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Linda" nameprefix="van de" lastname="Ree" gender="F" nation="NED" CLUB="De Ganze" birthdate="1963-10-26" />
    </RECORD>
    <RECORD swimtime="00:01:30.21">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rhenen" date="2023-03-18" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:03:12.07">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2023-01-07" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:00:33.64">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:01:19.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:03:08.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Margriet" nameprefix="" lastname="Grove-Lingeman" gender="F" nation="NED" CLUB="Triton" birthdate="1962-02-05" />
    </RECORD>
    <RECORD swimtime="00:01:16.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:02:45.80">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Rhenen" date="2023-03-18" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:06:04.89">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Almere-Poort" date="2023-03-12" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:28.88">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Glasgow" date="2023-04-22" nation="GBR" />
     <ATHLETE firstname="Dawn" nameprefix="" lastname="Kissack" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:05.34">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Castellon" date="2021-04-09" nation="ESP" />
     <ATHLETE firstname="Carmen" nameprefix="" lastname="Navarro" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:24.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Madrid" date="2022-01-15" nation="ESP" />
     <ATHLETE firstname="Carmen" nameprefix="" lastname="Navarro" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:05:09.41">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Palma de Mallorca" date="2022-04-23" nation="ESP" />
     <ATHLETE firstname="Barbara" nameprefix="" lastname="Gellrich" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:10:34.62">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-29" nation="GBR" />
     <ATHLETE firstname="Suzanne" nameprefix="" lastname="Noble" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:20:19.11">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-27" nation="GBR" />
     <ATHLETE firstname="Suzanne" nameprefix="" lastname="Noble" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:33.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <ATHLETE firstname="Julie" nameprefix="" lastname="Hoyle" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:13.93">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2022-10-28" nation="GBR" />
     <ATHLETE firstname="Julie" nameprefix="" lastname="Hoyle" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:38.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Glasgow" date="2022-04-08" nation="GBR" />
     <ATHLETE firstname="Julie" nameprefix="" lastname="Hoyle" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:37.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Castellon" date="2023-02-17" nation="ESP" />
     <ATHLETE firstname="Ute" nameprefix="" lastname="Hasse" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:21.14">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Trevisio" date="2022-04-14" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:03:00.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Molinela" date="2022-04-25" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:32.04">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Pontevedra" date="2022-01-15" nation="ESP" />
     <ATHLETE firstname="Carmen" nameprefix="" lastname="Navarro" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:11.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Castellon" date="2021-05-11" nation="ESP" />
     <ATHLETE firstname="Carmen" nameprefix="" lastname="Navarro" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:46.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Glasgow" date="2021-09-11" nation="SCO" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Pearson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:16.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Carlisle" date="2020-02-20" nation="GBR" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Pearson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:44.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Carlisle" date="2023-02-11" nation="GBR" />
     <ATHLETE firstname="Julie" nameprefix="" lastname="Hoyle" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:05:57.07">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Glasgow" date="2022-04-08" nation="GBR" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Pearson" gender="F" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:28.50">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-05-26" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:02.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-10-13" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:02:15.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-10-13" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:04:48.80">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-03-19" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:09:55.61">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-03-18" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:18:52.68">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-01-21" nation="CAN" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:00:32.91">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-04-23" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:12.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-10-13" nation="" />
     <ATHLETE firstname="Bonnie" nameprefix="" lastname="Bilich" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:34.31">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-04-24" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:37.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-05-26" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:20.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-05-26" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:02:57.05">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-05-26" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:00:31.24">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-07-12" nation="" />
     <ATHLETE firstname="Traci" nameprefix="" lastname="Granger" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:10.97">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-04-23" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:41.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2011-12-03" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:12.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-04-24" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:36.81">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-10-13" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:05:37.15">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-03-27" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:30.73">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2021-11-14" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:01:08.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2021-11-14" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:02:34.02">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-20" nation="POR" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:05:35.77">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:11:24.77">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:21:47.72">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-23" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:00:38.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:01:20.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:02:56.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:00:43.66">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Steenwijk" date="2019-09-14" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:01:33.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:03:21.44">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:00:35.82">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Steenwijk" date="2022-04-02" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:01:27.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:03:50.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2020-01-04" nation="NED" />
     <ATHLETE firstname="Margriet" nameprefix="" lastname="Pasma" gender="F" nation="NED" CLUB="TriVia" birthdate="1955-06-28" />
    </RECORD>
    <RECORD swimtime="00:01:20.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Funchal" date="2023-11-19" nation="POR" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:03:03.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Papendrecht" date="2023-01-07" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:06:54.20">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Almere-Poort" date="2023-03-12" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:29.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-28" nation="GBR" />
     <ATHLETE firstname="Alyson" nameprefix="" lastname="Fordham" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:07.07">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-29" nation="GBR" />
     <ATHLETE firstname="Alyson" nameprefix="" lastname="Fordham" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:33.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2022-10-28" nation="GBR" />
     <ATHLETE firstname="Alyson" nameprefix="" lastname="Fordham" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:05:19.64">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2020-01-26" nation="ITA" />
     <ATHLETE firstname="Cristina" nameprefix="" lastname="Tarantino" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:10:57.88">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2020-02-15" nation="ITA" />
     <ATHLETE firstname="Cristina" nameprefix="" lastname="Tarantino" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:20:51.88">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2020-02-08" nation="ITA" />
     <ATHLETE firstname="Cristina" nameprefix="" lastname="Tarantino" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:36.58">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="V�xj�" date="2010-03-21" nation="SWE" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:01:18.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2023-10-28" nation="GBR" />
     <ATHLETE firstname="Alyson" nameprefix="" lastname="Fordham" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:53.87">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Barnet Copthall" date="2023-07-09" nation="GBR" />
     <ATHLETE firstname="Alyson" nameprefix="" lastname="Fordham" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:38.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Essen" date="2021-11-28" nation="GER" />
     <ATHLETE firstname="Dagmar" nameprefix="" lastname="Frese" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:27.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2023-10-27" nation="GBR" />
     <ATHLETE firstname="Amanda" nameprefix="" lastname="Heath" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:07.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Crawley" date="2022-10-01" nation="GBR" />
     <ATHLETE firstname="Amanda" nameprefix="" lastname="Heath" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:35.38">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rostock" date="2019-05-18" nation="GER" />
     <ATHLETE firstname="Angela" nameprefix="" lastname="Zingler" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:23.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Wuppertal" date="2011-11-05" nation="GER" />
     <ATHLETE firstname="Brigitte" nameprefix="" lastname="Merten" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:06.07">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Palma de Mallorca" date="2024-01-14" nation="ESP" />
     <ATHLETE firstname="Ramona" nameprefix="" lastname="Guillen Munoz" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:19.69">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2023-10-29" nation="GBR" />
     <ATHLETE firstname="Alyson" nameprefix="" lastname="Fordham" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:57.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Palma de Mallorca" date="2024-01-13" nation="ESP" />
     <ATHLETE firstname="Ramona" nameprefix="" lastname="Guillen Munoz" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:06:21.67">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2022-10-28" nation="GBR" />
     <ATHLETE firstname="Amanda" nameprefix="" lastname="Heath" gender="F" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:29.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-11-19" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:04.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-01-12" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:23.26">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-11-18" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:02.08">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-09-24" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:10:34.67">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-01-30" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:20:05.72">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-01-28" nation="USA" />
     <ATHLETE firstname="Suzanne" nameprefix="" lastname="Heim-Bowen" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:33.41">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-09-22" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:13.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-01-12" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:42.87">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-12-01" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:38.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-11-28" nation="" />
     <ATHLETE firstname="Dagmar" nameprefix="" lastname="Frese" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:27.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-10-27" nation="" />
     <ATHLETE firstname="Amanda" nameprefix="" lastname="Heath" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:07.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-10-01" nation="" />
     <ATHLETE firstname="Amanda" nameprefix="" lastname="Heath" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:32.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-11-23" nation="" />
     <ATHLETE firstname="Penny" nameprefix="" lastname="Noyes" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:13.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-08-12" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:45.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2016-09-18" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:15.65">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-11-23" nation="" />
     <ATHLETE firstname="Penny" nameprefix="" lastname="Noyes" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:46.04">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-06-12" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:55.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-09-18" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:32.47">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:01:13.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:02:41.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:06:00.79">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:12:05.88">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:25:47.07">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-23" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:00:44.39">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:01:37.24">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:03:27.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kampen" date="2023-09-30" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:00:45.56">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Bea" nameprefix="" lastname="Swijnenberg" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1949-02-03" />
    </RECORD>
    <RECORD swimtime="00:01:41.53">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:03:46.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <ATHLETE firstname="Bea" nameprefix="" lastname="Swijnenberg" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1949-02-03" />
    </RECORD>
    <RECORD swimtime="00:00:38.89">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:01:40.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:04:36.06">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2020-01-04" nation="NED" />
     <ATHLETE firstname="Antoinette" nameprefix="" lastname="Gilding-Tussaud" gender="F" nation="NED" CLUB="WS Twente" birthdate="1950-05-19" />
    </RECORD>
    <RECORD swimtime="00:01:30.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Oss" date="2022-09-25" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:03:27.73">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:08:42.71">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2020-02-08" nation="NED" />
     <ATHLETE firstname="Antoinette" nameprefix="" lastname="Gilding-Tussaud" gender="F" nation="NED" CLUB="WS Twente" birthdate="1950-05-19" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:32.47">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:13.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:41.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:06:00.34">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Barnet" date="2003-09-28" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:12:05.88">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:23:54.74">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2004-11-28" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:37.50">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Stockholm" date="2015-03-21" nation="SWE" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:01:22.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Stockholm" date="2015-03-22" nation="SWE" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:03:05.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="London" date="2015-07-12" nation="GBR" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:00:42.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2023-04-22" nation="ITA" />
     <ATHLETE firstname="Carole Wendy" nameprefix="" lastname="Smith" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:34.86">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2014-10-25" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:28.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2014-10-24" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:36.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rennes" date="2015-03-25" nation="FRA" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:24.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Epinal" date="2016-01-30" nation="GBR" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:26.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Saransk" date="2018-11-17" nation="RUS" />
     <ATHLETE firstname="Kira" nameprefix="" lastname="Makarova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:23.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Palma de Mallorca" date="2016-04-02" nation="ESP" />
     <ATHLETE firstname="Brigitte" nameprefix="" lastname="Merten" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:11.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gau Algesheim" date="2016-01-17" nation="GER" />
     <ATHLETE firstname="Brigitte" nameprefix="" lastname="Merten" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:06:47.91">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gau Algesheim" date="2016-01-17" nation="GER" />
     <ATHLETE firstname="Brigitte" nameprefix="" lastname="Merten" gender="F" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:30.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-12-03" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:06.61">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-12-02" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:27.89">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-10-09" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:18.26">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-02-26" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:11:54.61">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2020-01-18" nation="" />
     <ATHLETE firstname="Cecilia" nameprefix="" lastname="Mccloskey" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:22:06.78">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2020-01-18" nation="" />
     <ATHLETE firstname="Cecilia" nameprefix="" lastname="Mccloskey" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:33.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-12-04" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:13.66">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-12-03" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:47.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-17" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:42.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-04-22" nation="" />
     <ATHLETE firstname="Carole Wendy" nameprefix="" lastname="Smith" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:33.92">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2015-04-12" nation="" />
     <ATHLETE firstname="Nobuko" nameprefix="" lastname="Yasuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:24.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-01-21" nation="" />
     <ATHLETE firstname="Nobuko" nameprefix="" lastname="Yasuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:34.14">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-02-25" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:15.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-10-17" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:57.32">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-10-07" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:18.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-12-04" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:52.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-10-16" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:07.14">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-10-06" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:36.72">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Oostburg" date="2021-10-30" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:01:27.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:03:13.82">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:07:13.95">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vlaardingen" date="2010-01-23" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:15:08.79">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2012-01-27" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:32:45.33">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-19" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:00:50.73">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Hoogerheide" date="2010-02-07" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:56.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2011-12-10" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:04:04.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Deurne" date="2010-04-18" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:00:48.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Funchal" date="2023-11-20" nation="POR" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:01:53.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Gemeentelijk zwembad Kapellen" date="2023-01-28" nation="BEL" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:04:02.10">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2023-01-07" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:00:57.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Oostburg" date="2021-10-30" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:03:12.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2011-01-23" nation="NED" />
     <ATHLETE firstname="Annie" nameprefix="de" lastname="Vos" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1934-01-10" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:44.57">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Oostburg" date="2021-10-30" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:03:49.82">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Oostburg" date="2021-10-30" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:10:46.66">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2011-01-23" nation="NED" />
     <ATHLETE firstname="Annie" nameprefix="de" lastname="Vos" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1934-01-10" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:34.58">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rostock" date="2015-06-20" nation="GER" />
     <ATHLETE firstname="Christel" nameprefix="" lastname="Schulz" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:18.59">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Guernsey" date="2006-03-25" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:57.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heron" date="2006-04-02" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:06:09.40">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2006-10-28" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:12:42.75">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2006-07-08" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:24:04.75">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Barnet" date="2006-11-26" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:40.74">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Lund" date="2018-02-17" nation="DEN" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:01:29.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Jarfalla" date="2020-01-11" nation="SWE" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:03:20.26">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Brondby" date="2018-03-11" nation="DEN" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:00:45.37">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2019-10-27" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:38.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Gelsenkirchen" date="2015-11-07" nation="GER" />
     <ATHLETE firstname="Luise" nameprefix="" lastname="Kn�pfle" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:36.11">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Gelsenkirchen" date="2015-11-07" nation="GER" />
     <ATHLETE firstname="Luise" nameprefix="" lastname="Kn�pfle" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:38.17">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Dunkerque" date="2019-03-08" nation="FRA" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:30.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Dunkerque" date="2019-03-09" nation="FRA" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:57.33">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Salzburg" date="2005-05-21" nation="AUT" />
     <ATHLETE firstname="Sylvia" nameprefix="" lastname="Neuhauser" gender="F" nation="AUT" />
    </RECORD>
    <RECORD swimtime="00:01:28.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="St. Petersburg" date="2022-01-09" nation="RUS" />
     <ATHLETE firstname="Kira" nameprefix="" lastname="Makarova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:03:28.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Berlin" date="2022-08-17" nation="GER" />
     <ATHLETE firstname="Brigitte" nameprefix="" lastname="Merten" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:07:34.39">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="London" date="2006-07-09" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:34.04">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-10-15" nation="" />
     <ATHLETE firstname="Diann" nameprefix="" lastname="Uustal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:15.87">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-17" nation="" />
     <ATHLETE firstname="Diann" nameprefix="" lastname="Uustal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:51.46">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-10-14" nation="" />
     <ATHLETE firstname="Diann" nameprefix="" lastname="Uustal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:08.74">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-04-19" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:12:25.61">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-05-12" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:24:04.75">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Barnet" date="2006-11-26" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:39.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-07-21" nation="" />
     <ATHLETE firstname="Clary" nameprefix="" lastname="Munns" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:26.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-10-15" nation="" />
     <ATHLETE firstname="Diann" nameprefix="" lastname="Uustal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:10.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-17" nation="" />
     <ATHLETE firstname="Diann" nameprefix="" lastname="Uustal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:43.79">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-02-14" nation="" />
     <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:36.48">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-03-21" nation="" />
     <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:33.03">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-04-17" nation="" />
     <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:38.17">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-08-03" nation="" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:30.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-09-03" nation="" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:34.50">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-05-25" nation="" />
     <ATHLETE firstname="Clary" nameprefix="" lastname="Munns" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:27.96">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-05-25" nation="" />
     <ATHLETE firstname="Clary" nameprefix="" lastname="Munns" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:03:15.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-11-13" nation="" />
     <ATHLETE firstname="Kira" nameprefix="" lastname="Makarova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:07:11.33">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2013-05-11" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:42.16">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-21" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:35.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:03:37.54">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2015-01-23" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:08:02.96">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:16:44.79">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-21" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:32:32.27">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-24" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:00:55.58">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:02:00.97">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Alphen" date="2018-09-15" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:04:19.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Roermond" date="2016-11-06" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:04.25">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roermond" date="2016-11-06" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:02:30.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Terneuzen" date="2009-09-10" nation="NED" />
     <ATHLETE firstname="Anneke" nameprefix="" lastname="Logtenberg" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1929-10-31" />
    </RECORD>
    <RECORD swimtime="00:05:27.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Breda" date="2001-01-28" nation="NED" />
     <ATHLETE firstname="Gr�" nameprefix="" lastname="Sch�nberger-de Hooge" gender="F" nation="NED" CLUB="ZPB H&amp;L Productions" birthdate="1921-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:03.78">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Mol" date="2019-10-05" nation="BEL" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:02:28.76">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:14.61">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Veldhoven" date="2015-02-08" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:37.67">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Guildford" date="2011-06-25" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:24.44">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Guildford" date="2011-06-25" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:01.61">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Guildford" date="2011-06-25" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:06:34.92">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Guernsey" date="2011-04-08" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:12:49.43">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Jersey" date="2011-06-11" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:25:45.37">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Jersey" date="2011-06-11" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:43.72">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Copenhagen" date="2023-10-01" nation="DEN" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:01:35.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Copenhagen" date="2023-09-30" nation="DEN" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:03:42.88">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="London" date="2011-07-17" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:47.20">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Portsmouth" date="2023-06-24" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:42.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Portsmouth" date="2023-06-24" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:53.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2023-10-29" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:45.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Guernsey" date="2011-04-09" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:59.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="London" date="2011-07-17" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:05:20.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Clermont" date="2010-03-11" nation="FRA" />
     <ATHLETE firstname="Yvette" nameprefix="" lastname="Kaplan Bader" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:42.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Guernsey" date="2011-04-10" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:43.73">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Jersey" date="2011-06-11" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:07.34">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="London" date="2011-07-17" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:36.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-05-20" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:21.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-05-20" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:00.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-10-02" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:06:23.17">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-10-20" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:12:49.43">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-11-06" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:25:45.37">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-06-11" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:43.76">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-05-15" nation="" />
     <ATHLETE firstname="Satoko" nameprefix="" lastname="Takeuji" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:35.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-09-30" nation="" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:03:32.48">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-03-19" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Yoshida" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:46.48">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2015-03-08" nation="" />
     <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:42.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-06-24" nation="" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:53.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-10-28" nation="" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:45.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Guernsey" date="2011-04-09" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:50.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2012-04-01" nation="" />
     <ATHLETE firstname="Judie" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:04:10.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2012-03-31" nation="" />
     <ATHLETE firstname="Judie" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:38.45">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-01-20" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:43.73">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2011-06-11" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:04.67">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2012-03-30" nation="" />
     <ATHLETE firstname="Judie" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:48.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-21" nation="POR" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:49.72">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:04:01.16">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:08:44.87">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roermond" date="2023-09-24" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:17:47.07">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Veldhoven" date="2023-06-04" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:35:58.75">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-16" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:00:59.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:02:16.32">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Funchal" date="2023-11-21" nation="POR" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:06:57.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Geel" date="2013-06-08" nation="BEL" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:01:07.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Leiden" date="2024-01-21" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:02:35.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Maastricht" date="2023-12-28" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:06:40.21">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2011-02-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:01:10.53">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Veldhoven" date="2023-06-04" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:02:40.62">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Maastricht" date="2023-12-29" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:17.83">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Etten-Leur" date="2023-11-05" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:37.75">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Guernsey" date="2016-04-17" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:28.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Guildford" date="2016-06-25" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:12.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Guildford" date="2016-06-25" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:06:57.06">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Guernsey" date="2016-04-15" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:15:33.71">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gau-Algesheim" date="2023-01-14" nation="GER" />
     <ATHLETE firstname="Helga" nameprefix="" lastname="Reich" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:28:02.25">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2016-11-27" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:47.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Szazhalombatta" date="2019-02-24" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:01:44.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Szazhalombatta" date="2019-02-23" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:03:48.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Szazhalombatta" date="2019-02-24" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:00:52.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2016-01-23" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:01:56.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:04:17.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Nijlen" date="2016-03-19" nation="BEL" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:00:51.79">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Szazhalombatta" date="2020-02-15" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:01.30">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Szazhalombatta" date="2020-02-16" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:06:04.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Colmar" date="2014-02-02" nation="FRA" />
     <ATHLETE firstname="Yvette" nameprefix="" lastname="Kaplan Bader" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:47.02">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Inverness" date="2016-08-20" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:57.27">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Szazhalombatta" date="2019-02-23" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:12:39.03">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Erstein " date="2014-05-01" nation="FRA" />
     <ATHLETE firstname="Yvette" nameprefix="" lastname="Kaplan Bader" gender="F" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:38.75">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-04-17" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:27.19">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-04-08" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:12.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-06-25" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:06:57.06">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-04-15" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:14:24.83">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-09-16" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:28:02.25">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-11-27" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:45.54">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-05-28" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:43.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-07-02" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:48.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-02-24" nation="" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:00:52.17">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2016-01-23" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:01:56.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:04:17.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-03-19" nation="" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:00:51.40">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-03-25" nation="" />
     <ATHLETE firstname="Judie" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:02:02.59">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-05-12" nation="" />
     <ATHLETE firstname="Judie" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:04:40.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-03-25" nation="" />
     <ATHLETE firstname="Judie" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:47.02">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-08-20" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:57.27">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-02-23" nation="" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:08:42.45">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-03-24" nation="" />
     <ATHLETE firstname="Judie" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:01:16.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2016-01-09" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:06.83">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:07:15.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Andel" date="2016-03-13" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:27.72">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwolle" date="2016-01-09" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:27.52">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2017-12-02" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:07:19.81">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2017-12-02" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:01:37.78">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:29.73">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:08:40.58">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-12-03" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:00:45.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2021-10-30" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:44.21">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2021-10-29" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:54.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2021-10-30" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:48.34">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2021-11-28" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:17:58.34">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:33:41.77">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2021-11-28" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:04.17">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eskilstuna" date="2017-03-26" nation="SWE" />
     <ATHLETE firstname="Kerstin" nameprefix="" lastname="Gj�res" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:02:01.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2021-10-31" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:05:02.82">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2006-10-28" nation="GBR" />
     <ATHLETE firstname="Willy" nameprefix="van" lastname="Rysel" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:58.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Embourg" date="2023-03-19" nation="BEL" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:02:09.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Embourg" date="2023-03-18" nation="BEL" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:04:44.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Embourg" date="2023-03-18" nation="BEL" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:01:34.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Isle of Wight" date="2003-02-22" nation="GBR" />
     <ATHLETE firstname="Dorothy" nameprefix="" lastname="Weston" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:21.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Guernsey" date="2003-04-06" nation="GBR" />
     <ATHLETE firstname="Dorothy" nameprefix="" lastname="Weston" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="00:02:09.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:00:45.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-30" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:44.21">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-29" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:52.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-02" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:48.34">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-11-28" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:17:58.34">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-11-28" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:33:41.77">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-11-28" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:55.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-02" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:01.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-31" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:04:24.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-10-15" nation="" />
     <ATHLETE firstname="Betty" nameprefix="" lastname="Lorenzi" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:59.04">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2023-11-26" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:02:13.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2023-11-26" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:05:15.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Chartres" date="2013-03-07" nation="FRA" />
     <ATHLETE firstname="Olga" nameprefix="" lastname="Kokorina" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:02.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-12-18" nation="" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:02:28.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-04-24" nation="" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:05:33.79">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-11-06" nation="" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:02:09.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-10-29" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:04:50.01">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-04-24" nation="" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:10:29.18">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-11-06" nation="" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:01:25.93">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2022-09-24" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:43.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Oostburg" date="2021-10-30" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:08:26.16">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:40.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:46.31">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Etten-Leur" date="2022-11-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:08:07.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Etten-Leur" date="2022-11-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:02:02.87">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:04:43.59">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Oostburg" date="2021-10-30" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:09:48.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Oostburg" date="2021-10-30" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:01:07.27">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kaerepere" date="2017-02-04" nation="EST" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Kutti" gender="F" nation="EST" />
    </RECORD>
    <RECORD swimtime="00:03:43.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Caen" date="2016-03-06" nation="FRA" />
     <ATHLETE firstname="Michele" nameprefix="" lastname="Guillais" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:08:26.16">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:19:24.06">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Palma de Mallorca" date="2006-04-23" nation="ESP" />
     <ATHLETE firstname="Rosa" nameprefix="" lastname="Sellares" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="00:01:12.24">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kaerepere" date="2017-02-04" nation="EST" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Kutti" gender="F" nation="EST" />
    </RECORD>
    <RECORD swimtime="00:02:53.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Tallinn" date="2017-04-09" nation="EST" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Kutti" gender="F" nation="EST" />
    </RECORD>
    <RECORD swimtime="00:08:07.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Etten-Leur" date="2022-11-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:26.91">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Hannover" date="2016-11-26" nation="GER" />
     <ATHLETE firstname="Ingeborg" nameprefix="" lastname="Fritze" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:43.54">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Oostburg" date="2021-10-30" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:09:48.06">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Oostburg" date="2021-10-30" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:01:00.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-04-22" nation="" />
     <ATHLETE firstname="Elizabeth" nameprefix="" lastname="Wallis" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:02:16.63">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-12-01" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:56.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-01-12" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:10:08.44">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-12-03" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:20:57.02">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-11-06" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:42:34.14">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-10-06" nation="" />
     <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:12.24">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-02-04" nation="" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Kutti" gender="F" nation="EST" />
    </RECORD>
    <RECORD swimtime="00:02:42.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-04-27" nation="" />
     <ATHLETE firstname="Kalis" nameprefix="" lastname="Rasmussen" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:05:42.83">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-04-28" nation="" />
     <ATHLETE firstname="Kalis" nameprefix="" lastname="Rasmussen" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:32.51">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-04-28" nation="" />
     <ATHLETE firstname="Kalis" nameprefix="" lastname="Rasmussen" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:03:33.94">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-04-28" nation="" />
     <ATHLETE firstname="Kalis" nameprefix="" lastname="Rasmussen" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:07:22.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-04-28" nation="" />
     <ATHLETE firstname="Kalis" nameprefix="" lastname="Rasmussen" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:02:12.78">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-12-02" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="00:03:32.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-09-25" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:32.59">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-10-12" nation="" />
     <ATHLETE firstname="Charlotte" nameprefix="" lastname="Sanddal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="00:03:53.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Barcelona" date="2010-01-09" nation="ESP" />
     <ATHLETE firstname="Rosa" nameprefix="" lastname="Sellares" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="00:01:15.61">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-03" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:30.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-01-26" nation="" />
     <ATHLETE firstname="Mieko" nameprefix="" lastname="Nagaoka" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:07:27.89">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-01-25" nation="" />
     <ATHLETE firstname="Mieko" nameprefix="" lastname="Nagaoka" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:16:40.10">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-04-06" nation="" />
     <ATHLETE firstname="Mieko" nameprefix="" lastname="Nagaoka" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:36:51.23">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-05-11" nation="" />
     <ATHLETE firstname="Mieko" nameprefix="" lastname="Nagaoka" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="01:15:54.39">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-04-04" nation="" />
     <ATHLETE firstname="Mieko" nameprefix="" lastname="Nagaoka" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:29.22">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-03" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:55.51">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-03" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:22.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-03" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="00:06:02.24">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-10-06" nation="" />
     <ATHLETE firstname="Charlotte" nameprefix="" lastname="Sanddal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:12:48.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-10-05" nation="" />
     <ATHLETE firstname="Charlotte" nameprefix="" lastname="Sanddal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="00:05:01.09">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-10-06" nation="" />
     <ATHLETE firstname="Charlotte" nameprefix="" lastname="Sanddal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="20" agemax="24" />
   <RECORDS>
    <RECORD swimtime="00:00:22.76">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="startlimiet" nameprefix="" lastname="" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:50.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="startlimiet" nameprefix="" lastname="" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:52.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2015-02-21" nation="NED" />
     <ATHLETE firstname="Kevin" nameprefix="" lastname="Eltink" gender="M" nation="NED" CLUB="DWK" birthdate="1991-10-29" />
    </RECORD>
    <RECORD swimtime="00:04:03.40">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2014-12-22" nation="NED" />
     <ATHLETE firstname="Fabian" nameprefix="" lastname="Beimin" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1991-06-08" />
    </RECORD>
    <RECORD swimtime="00:08:19.90">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2014-12-22" nation="NED" />
     <ATHLETE firstname="Fabian" nameprefix="" lastname="Beimin" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1991-06-08" />
    </RECORD>
    <RECORD swimtime="00:15:59.90">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2014-12-22" nation="NED" />
     <ATHLETE firstname="Fabian" nameprefix="" lastname="Beimin" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1991-06-08" />
    </RECORD>
    <RECORD swimtime="00:00:26.33">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Vlissingen" date="2009-01-25" nation="NED" />
     <ATHLETE firstname="Merijn" nameprefix="" lastname="Ellenkamp" gender="M" nation="NED" CLUB="DWK" birthdate="1985-06-30" />
    </RECORD>
    <RECORD swimtime="00:00:57.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Vlissingen" date="2009-01-24" nation="NED" />
     <ATHLETE firstname="Merijn" nameprefix="" lastname="Ellenkamp" gender="M" nation="NED" CLUB="DWK" birthdate="1985-06-30" />
    </RECORD>
    <RECORD swimtime="00:02:04.41">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Terneuzen" date="2012-01-27" nation="NED" />
     <ATHLETE firstname="Jos" nameprefix="de" lastname="Graaf" gender="M" nation="NED" CLUB="PSV" birthdate="1991-08-31" />
    </RECORD>
    <RECORD swimtime="00:00:28.67">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2023-11-26" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="" lastname="Peters" gender="M" nation="NED" CLUB="Nuenen" birthdate="1999-02-24" />
    </RECORD>
    <RECORD swimtime="00:01:03.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <ATHLETE firstname="Jordan" nameprefix="" lastname="Kraaijenhof" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1993-07-16" />
    </RECORD>
    <RECORD swimtime="00:02:19.77">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Jordan" nameprefix="" lastname="Kraaijenhof" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1993-07-16" />
    </RECORD>
    <RECORD swimtime="00:00:24.17">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Verhoeven" gender="M" nation="NED" CLUB="Albion WSS (SG)" birthdate="1997-04-18" />
    </RECORD>
    <RECORD swimtime="00:00:55.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Verhoeven" gender="M" nation="NED" CLUB="Albion WSS (SG)" birthdate="1997-04-18" />
    </RECORD>
    <RECORD swimtime="00:02:07.31">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2014-01-25" nation="NED" />
     <ATHLETE firstname="Kevin" nameprefix="" lastname="Eltink" gender="M" nation="NED" CLUB="DWK" birthdate="1991-10-29" />
    </RECORD>
    <RECORD swimtime="00:00:56.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="startlimiet" nameprefix="" lastname="" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:06.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2015-01-23" nation="NED" />
     <ATHLETE firstname="Kevin" nameprefix="" lastname="Eltink" gender="M" nation="NED" CLUB="DWK" birthdate="1991-10-29" />
    </RECORD>
    <RECORD swimtime="00:04:33.61">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2015-01-24" nation="NED" />
     <ATHLETE firstname="Kevin" nameprefix="" lastname="Eltink" gender="M" nation="NED" CLUB="DWK" birthdate="1991-10-29" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:22.38">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:00:50.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2008-12-13" nation="NED" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Oosting" gender="M" nation="NED" CLUB="PSV" birthdate="1981-04-01" />
    </RECORD>
    <RECORD swimtime="00:01:52.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-23" nation="NED" />
     <ATHLETE firstname="Kevin" nameprefix="" lastname="Eltink" gender="M" nation="NED" CLUB="DWK" birthdate="1991-10-29" />
    </RECORD>
    <RECORD swimtime="00:04:06.04">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2012-01-28" nation="NED" />
     <ATHLETE firstname="Raymond" nameprefix="van der" lastname="Merwe" gender="M" nation="NED" CLUB="WVZ" birthdate="1986-11-19" />
    </RECORD>
    <RECORD swimtime="00:08:42.72">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vlaardingen" date="2010-01-24" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:16:34.60">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2011-01-23" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:00:25.25">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Albion WSS (SG)" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:00:54.62">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Albion WSS (SG)" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:02:04.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Terneuzen" date="2012-01-27" nation="NED" />
     <ATHLETE firstname="Raymond" nameprefix="van der" lastname="Merwe" gender="M" nation="NED" CLUB="WVZ" birthdate="1986-11-19" />
    </RECORD>
    <RECORD swimtime="00:00:28.52">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Dominique" nameprefix="" lastname="Sikkema" gender="M" nation="NED" CLUB="TriVia" birthdate="1995-01-24" />
    </RECORD>
    <RECORD swimtime="00:01:03.31">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" CLUB="De Kempvis" birthdate="1993-08-07" />
    </RECORD>
    <RECORD swimtime="00:02:22.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2016-01-24" nation="NED" />
     <ATHLETE firstname="Kevin" nameprefix="" lastname="Eltink" gender="M" nation="NED" CLUB="DWK" birthdate="1991-10-29" />
    </RECORD>
    <RECORD swimtime="00:00:24.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:00:55.22">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:02:05.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Maastricht" date="2017-01-20" nation="NED" />
     <ATHLETE firstname="Kevin" nameprefix="" lastname="Eltink" gender="M" nation="NED" CLUB="DWK" birthdate="1991-10-29" />
    </RECORD>
    <RECORD swimtime="00:00:55.31">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Albion WSS (SG)" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:02:05.88">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <ATHLETE firstname="Kevin" nameprefix="" lastname="Eltink" gender="M" nation="NED" CLUB="DWK" birthdate="1991-10-29" />
    </RECORD>
    <RECORD swimtime="00:04:28.38">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Terneuzen" date="2012-01-29" nation="NED" />
     <ATHLETE firstname="Raymond" nameprefix="van der" lastname="Merwe" gender="M" nation="NED" CLUB="WVZ" birthdate="1986-11-19" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:21.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Jyv�skyl�" date="2014-09-13" nation="FIN" />
     <ATHLETE firstname="Ari-Pekka" nameprefix="" lastname="Liukkonen" gender="M" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:00:48.58">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Hildesheim" date="2005-11-19" nation="GER" />
     <ATHLETE firstname="Stephan" nameprefix="" lastname="Kunzelmann" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:49.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Malaga" date="2018-02-04" nation="ESP" />
     <ATHLETE firstname="David" nameprefix="" lastname="Alcolado" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:03:51.56">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Newport" date="2023-12-02" nation="GBR" />
     <ATHLETE firstname="William" nameprefix="" lastname="Ryley" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:13.81">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2003-10-24" nation="GBR" />
     <ATHLETE firstname="Greg" nameprefix="" lastname="Orphanides" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:15:29.68">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2003-10-24" nation="GBR" />
     <ATHLETE firstname="Greg" nameprefix="" lastname="Orphanides" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:23.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Tallin" date="2020-12-02" nation="EST" />
     <ATHLETE firstname="Ralf" nameprefix="" lastname="Tribuntsov" gender="M" nation="EST" />
    </RECORD>
    <RECORD swimtime="00:00:54.05">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Torino" date="2023-12-09" nation="ITA" />
     <ATHLETE firstname="Emanuel" nameprefix="" lastname="Turchi" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:56.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kiel" date="2006-12-16" nation="GER" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Herbst" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:26.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2017-10-29" nation="GBR" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Palmer" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:59.23">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2017-10-28" nation="GBR" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Palmer" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:11.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2017-10-27" nation="GBR" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Palmer" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:23.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="2021-10-31" nation="GBR" />
     <ATHLETE firstname="Adam" nameprefix="" lastname="Barrett" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:51.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="2021-10-29" nation="GBR" />
     <ATHLETE firstname="Adam" nameprefix="" lastname="Barrett" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:59.74">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Guildford" date="2008-09-20" nation="GBR" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Lewis" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:55.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Tallinn" date="2017-04-08" nation="EST" />
     <ATHLETE firstname="Martin" nameprefix="" lastname="Liivamaegi" gender="M" nation="EST" />
    </RECORD>
    <RECORD swimtime="00:01:58.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2019-11-22" nation="RUS" />
     <ATHLETE firstname="Dmitri" nameprefix="" lastname="Gorbunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:04:19.10">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Newport" date="2023-12-03" nation="GBR" />
     <ATHLETE firstname="William" nameprefix="" lastname="Ryley" gender="M" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:21.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-11-20" nation="" />
     <ATHLETE firstname="Ryan" nameprefix="" lastname="Held" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:47.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-11-16" nation="" />
     <ATHLETE firstname="Cesar" nameprefix="" lastname="Cielo" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:44.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-11-03" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:52.83">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-12-09" nation="" />
     <ATHLETE firstname="Drew" nameprefix="" lastname="Modrov" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:07.91">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2001-04-12" nation="" />
     <ATHLETE firstname="Alexandre" nameprefix="" lastname="Angelotti" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:15:29.68">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2003-10-24" nation="GBR" />
     <ATHLETE firstname="Greg" nameprefix="" lastname="Orphanides" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:23.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-11-21" nation="" />
     <ATHLETE firstname="Ryan" nameprefix="" lastname="Held" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:52.05">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-01-14" nation="JPN" />
     <ATHLETE firstname="Ryota" nameprefix="" lastname="Maejima" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:56.01">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-01-15" nation="JPN" />
     <ATHLETE firstname="Ryota" nameprefix="" lastname="Maejima" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:26.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-10-29" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Palmer" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:58.14">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-11-28" nation="" />
     <ATHLETE firstname="Shotaro" nameprefix="" lastname="Shimazaki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:07.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-10-14" nation="" />
     <ATHLETE firstname="Josh" nameprefix="" lastname="Prenot" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:23.15">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-11-21" nation="" />
     <ATHLETE firstname="Ryan" nameprefix="" lastname="Held" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:51.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-10-29" nation="" />
     <ATHLETE firstname="Adam" nameprefix="" lastname="Barrett" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:53.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-03-21" nation="" />
     <ATHLETE firstname="Syun" nameprefix="" lastname="Watarai" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:52.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-11-21" nation="" />
     <ATHLETE firstname="Ryan" nameprefix="" lastname="Held" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:58.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2020-10-04" nation="" />
     <ATHLETE firstname="Ken" nameprefix="" lastname="Kuwayama" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:04:14.51">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-11-15" nation="" />
     <ATHLETE firstname="Ikumi" nameprefix="" lastname="Hasegawa" gender="M" nation="JPN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:22.82">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <ATHLETE firstname="Joan" nameprefix="" lastname="Kentrop" gender="M" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1985-12-01" />
    </RECORD>
    <RECORD swimtime="00:00:50.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-20" nation="NED" />
     <ATHLETE firstname="Joan" nameprefix="" lastname="Kentrop" gender="M" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1985-12-01" />
    </RECORD>
    <RECORD swimtime="00:01:56.59">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Lelystad" date="1997-03-15" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:10.97">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2015-01-24" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:08:41.47">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:16:38.05">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-19" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:00:26.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Racing Club" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:00:58.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Jesper" nameprefix="" lastname="Oranje" gender="M" nation="NED" CLUB="De Duck" birthdate="1992-05-15" />
    </RECORD>
    <RECORD swimtime="00:02:11.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Breda" date="1994-01-30" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:28.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Gavin" nameprefix="van der" lastname="Werf" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1993-10-11" />
    </RECORD>
    <RECORD swimtime="00:01:03.62">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Gavin" nameprefix="van der" lastname="Werf" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1993-10-11" />
    </RECORD>
    <RECORD swimtime="00:02:20.07">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Gavin" nameprefix="van der" lastname="Werf" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1993-10-11" />
    </RECORD>
    <RECORD swimtime="00:00:25.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Marc" nameprefix="" lastname="Kremer" gender="M" nation="NED" CLUB="ReVeLie Swim Team" birthdate="1990-10-25" />
    </RECORD>
    <RECORD swimtime="00:00:25.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Jesper" nameprefix="" lastname="Oranje" gender="M" nation="NED" CLUB="De Duck" birthdate="1992-05-15" />
    </RECORD>
    <RECORD swimtime="00:00:56.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Racing Club" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:02:11.59">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Maastricht" date="2017-01-20" nation="NED" />
     <ATHLETE firstname="Alex" nameprefix="" lastname="Schelvis" gender="M" nation="NED" CLUB="LINK" birthdate="1987-08-09" />
    </RECORD>
    <RECORD swimtime="00:00:57.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Racing Club" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:02:08.41">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Oss" date="1996-12-15" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:40.29">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Winterswijk" date="2002-05-04" nation="NED" />
     <ATHLETE firstname="Diederik" nameprefix="" lastname="Rouffaer" gender="M" nation="NED" CLUB="ZON/S&amp;S" birthdate="1972-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:21.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="St. Petersburg" date="2015-11-28" nation="RUS" />
     <ATHLETE firstname="Evgeni" nameprefix="" lastname="Lagunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:47.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="St. Petersburg" date="2015-11-27" nation="RUS" />
     <ATHLETE firstname="Evgeni" nameprefix="" lastname="Lagunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:46.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kiel" date="2011-12-17" nation="GER" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Herbst" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:48.54">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Copenhagen" date="2023-09-30" nation="DEN" />
     <ATHLETE firstname="Frans" nameprefix="" lastname="Johannessen" gender="M" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:08:06.56">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Copenhagen" date="2023-09-30" nation="DEN" />
     <ATHLETE firstname="Frans" nameprefix="" lastname="Johannessen" gender="M" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:16:00.22">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Onda" date="2017-05-13" nation="ESP" />
     <ATHLETE firstname="Rafael" nameprefix="" lastname="Cabanillas" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:24.68">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Saransk" date="2019-11-24" nation="RUS" />
     <ATHLETE firstname="Sergey" nameprefix="" lastname="Makov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:54.53">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Saransk" date="2019-11-22" nation="RUS" />
     <ATHLETE firstname="Sergey" nameprefix="" lastname="Makov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:56.68">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kiel" date="2008-12-20" nation="GER" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Herbst" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:27.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2015-11-27" nation="RUS" />
     <ATHLETE firstname="Sergei" nameprefix="" lastname="Geibel" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:59.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2015-11-28" nation="RUS" />
     <ATHLETE firstname="Sergei" nameprefix="" lastname="Geibel" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:11.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Saransk" date="2021-11-13" nation="RUS" />
     <ATHLETE firstname="Dmitryi" nameprefix="" lastname="Gobunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:22.87">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rostock" date="2009-05-16" nation="GER" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Rupprath" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:52.64">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Barcelona" date="2009-05-31" nation="ESP" />
     <ATHLETE firstname="Fernando" nameprefix="" lastname="Alaez" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:53.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Burevestnik" date="2017-11-25" nation="RUS" />
     <ATHLETE firstname="Nikolay" nameprefix="" lastname="Skvortsov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:54.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Olsztyn" date="2018-11-17" nation="POL" />
     <ATHLETE firstname="Pawel" nameprefix="" lastname="Korzeniowski" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:01:58.13">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Kiel" date="2008-12-20" nation="GER" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Herbst" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:24.21">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Copenhagen" date="2023-10-01" nation="DEN" />
     <ATHLETE firstname="Frans" nameprefix="" lastname="Johannessen" gender="M" nation="DEN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:21.53">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-12-05" nation="" />
     <ATHLETE firstname="F." nameprefix="" lastname="Rosa Messias" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:00:47.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-11-27" nation="" />
     <ATHLETE firstname="Evgeni" nameprefix="" lastname="Lagunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:46.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-09-27" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:48.54">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-09-30" nation="" />
     <ATHLETE firstname="Frans" nameprefix="" lastname="Johanessen" gender="M" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:08:06.56">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-09-30" nation="" />
     <ATHLETE firstname="Frans" nameprefix="" lastname="Johanessen" gender="M" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:15:30.92">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-01-26" nation="" />
     <ATHLETE firstname="Chad" nameprefix="la" lastname="Tourette" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:23.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-05-07" nation="" />
     <ATHLETE firstname="Nelson" nameprefix="" lastname="Silva jr." gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:00:52.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-02-13" nation="" />
     <ATHLETE firstname="Junichi" nameprefix="" lastname="Morita" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:53.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-03-12" nation="" />
     <ATHLETE firstname="Junichi" nameprefix="" lastname="Morita" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:26.72">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-05-05" nation="" />
     <ATHLETE firstname="Felipe" nameprefix="" lastname="Lima" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:00:59.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-11-28" nation="" />
     <ATHLETE firstname="Kohhei" nameprefix="" lastname="Tominaga" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:11.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-11-13" nation="" />
     <ATHLETE firstname="Dmitrii" nameprefix="" lastname="Gorbunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:22.87">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rostock" date="2009-05-16" nation="GER" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Rupprath" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:52.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-04-16" nation="" />
     <ATHLETE firstname="Ko" nameprefix="" lastname="Fukaya" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:53.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-11-25" nation="" />
     <ATHLETE firstname="Nikolay" nameprefix="" lastname="Skvortsov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:53.28">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-11-13" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:56.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-11-13" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:16.06">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-11-12" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:23.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Joan" nameprefix="" lastname="Kentrop" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1985-12-01" />
    </RECORD>
    <RECORD swimtime="00:00:51.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Joan" nameprefix="" lastname="Kentrop" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1985-12-01" />
    </RECORD>
    <RECORD swimtime="00:01:53.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Breda" date="1998-01-25" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:07.22">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="1998-01-10" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:08:46.81">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Apeldoorn" date="1999-02-20" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:16:56.13">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-24" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:00:27.22">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Joan" nameprefix="" lastname="Kentrop" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1985-12-01" />
    </RECORD>
    <RECORD swimtime="00:00:58.21">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1985-03-27" />
    </RECORD>
    <RECORD swimtime="00:02:09.92">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwolle" date="1999-01-09" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:27.93">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1985-03-27" />
    </RECORD>
    <RECORD swimtime="00:01:02.11">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1985-03-27" />
    </RECORD>
    <RECORD swimtime="00:02:16.82">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1985-03-27" />
    </RECORD>
    <RECORD swimtime="00:00:24.84">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1985-03-27" />
    </RECORD>
    <RECORD swimtime="00:00:56.44">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1985-03-27" />
    </RECORD>
    <RECORD swimtime="00:02:13.13">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zoetermeer" date="1996-01-20" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:00:56.07">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Rotterdam Swimming (SG)" birthdate="1985-03-27" />
    </RECORD>
    <RECORD swimtime="00:02:08.21">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Breda" date="1999-01-31" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:39.42">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Almere" date="1999-11-14" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:21.53">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2007-10-27" nation="GBR" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Foster" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:49.37">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Essen" date="2021-11-28" nation="GER" />
     <ATHLETE firstname="Stefano" nameprefix="" lastname="Razeto" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:51.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Bonn" date="2004-11-27" nation="GER" />
     <ATHLETE firstname="Jochen" nameprefix="" lastname="Bruha" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:58.46">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2017-04-23" nation="ITA" />
     <ATHLETE firstname="Nicola" nameprefix="" lastname="Nisato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:08:19.97">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Genova" date="2022-03-27" nation="ITA" />
     <ATHLETE firstname="Lorenzo" nameprefix="" lastname="Giovanni" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:15:58.12">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2022-12-04" nation="ITA" />
     <ATHLETE firstname="Giovanni" nameprefix="" lastname="Lorenzo" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:24.48">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Essen" date="2021-11-27" nation="GER" />
     <ATHLETE firstname="Stefano" nameprefix="" lastname="Razeto" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:54.59">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Castellon" date="2023-02-19" nation="ESP" />
     <ATHLETE firstname="Carlos" nameprefix="" lastname="Requeno Soler" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:01.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kiel" date="2013-12-14" nation="GER" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Herbst" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:27.32">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kazan" date="2016-11-18" nation="RUS" />
     <ATHLETE firstname="Sergei" nameprefix="" lastname="Geibel" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:00.61">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kazan" date="2016-11-19" nation="RUS" />
     <ATHLETE firstname="Sergei" nameprefix="" lastname="Geibel" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:16.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2004-10-30" nation="GBR" />
     <ATHLETE firstname="Nick" nameprefix="" lastname="Gillingham" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:23.63">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Essen" date="2021-11-27" nation="GER" />
     <ATHLETE firstname="Stefano" nameprefix="" lastname="Razeto" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:54.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2012-04-01" nation="ITA" />
     <ATHLETE firstname="Massimiliano" nameprefix="" lastname="Eroli" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:03.05">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2012-02-18" nation="ITA" />
     <ATHLETE firstname="Massimiliano" nameprefix="" lastname="Eroli" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:54.86">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Poznan" date="2022-12-17" nation="POL" />
     <ATHLETE firstname="Pawel" nameprefix="" lastname="Korzeniowski" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:02:05.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Lucca" date="2012-12-02" nation="ITA" />
     <ATHLETE firstname="Massimiliano" nameprefix="" lastname="Eroli" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:04:30.09">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Rundforbi" date="2015-03-08" nation="DEN" />
     <ATHLETE firstname="Claus" nameprefix="" lastname="Iversen" gender="M" nation="DEN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:21.53">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2007-10-27" nation="" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Foster" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:47.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-11-18" nation="" />
     <ATHLETE firstname="Roland" nameprefix="" lastname="Schoeman" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:48.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-12-02" nation="" />
     <ATHLETE firstname="Benjamin" nameprefix="" lastname="Hockin" gender="M" nation="PAR" />
    </RECORD>
    <RECORD swimtime="00:03:57.77">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2003-12-14" nation="" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Hochstein" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:16.19">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-12-06" nation="" />
     <ATHLETE firstname="Alex" nameprefix="" lastname="Kostich" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:15:41.78">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-01-28" nation="USA" />
     <ATHLETE firstname="Chad" nameprefix="la" lastname="Tourette" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:24.48">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-11-27" nation="" />
     <ATHLETE firstname="Stefano" nameprefix="" lastname="Razeto" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:54.59">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-02-19" nation="" />
     <ATHLETE firstname="Carlos" nameprefix="" lastname="Requeno Soler" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:00.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2002-12-08" nation="" />
     <ATHLETE firstname="Ron" nameprefix="" lastname="Karnaugh" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:26.66">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-11-17" nation="" />
     <ATHLETE firstname="Roland" nameprefix="" lastname="Schoeman" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:59.65">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-03-19" nation="" />
     <ATHLETE firstname="Ryo" nameprefix="" lastname="Kobayashi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:15.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2014-03-16" nation="" />
     <ATHLETE firstname="Kazuya" nameprefix="" lastname="Koike" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:23.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2018-11-18" nation="" />
     <ATHLETE firstname="Roland" nameprefix="" lastname="Schoeman" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:52.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2020-01-18" nation="" />
     <ATHLETE firstname="Takuya" nameprefix="" lastname="Hasegawa" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:00.01">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-05-28" nation="" />
     <ATHLETE firstname="Tatsuya" nameprefix="" lastname="Ito" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:54.86">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-12-17" nation="" />
     <ATHLETE firstname="Pawel" nameprefix="" lastname="Korzeniowski" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:01:59.85">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-10-27" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:19.79">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-10-26" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:23.74">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:00:51.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:01:58.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zuidbroek" date="2003-11-15" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:19.38">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1976-06-26" />
    </RECORD>
    <RECORD swimtime="00:08:53.53">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vlissingen" date="2008-03-02" nation="NED" />
     <ATHLETE firstname="Joost" nameprefix="" lastname="Kuijlaars" gender="M" nation="NED" CLUB="MNC Dordrecht" birthdate="1966-01-01" />
    </RECORD>
    <RECORD swimtime="00:17:29.80">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vlissingen" date="2006-02-19" nation="NED" />
     <ATHLETE firstname="Joost" nameprefix="" lastname="Kuijlaars" gender="M" nation="NED" CLUB="SBC2000" birthdate="1966-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:27.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" CLUB="De Lansingh" birthdate="1980-05-09" />
    </RECORD>
    <RECORD swimtime="00:00:59.94">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Grootebroek" date="2003-05-18" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:10.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Lelystad" date="2004-03-20" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:29.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2009-11-29" nation="NED" />
     <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" CLUB="PSV" birthdate="1968-10-13" />
    </RECORD>
    <RECORD swimtime="00:01:06.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Best" date="2009-09-27" nation="NED" />
     <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" CLUB="PSV" birthdate="1968-10-13" />
    </RECORD>
    <RECORD swimtime="00:02:27.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zuidbroek" date="2003-11-14" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:25.81">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:00:58.33">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:02:16.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zoetermeer" date="2000-04-01" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:00.19">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:02:12.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Emmeloord" date="2006-01-22" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:47.69">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Papendrecht" date="2016-01-24" nation="NED" />
     <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1976-06-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:22.39">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-21" nation="POR" />
     <ATHLETE firstname="Filippo" nameprefix="" lastname="Magnini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:48.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-23" nation="POR" />
     <ATHLETE firstname="Filippo" nameprefix="" lastname="Magnini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:49.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Milano" date="2023-12-17" nation="ITA" />
     <ATHLETE firstname="Filippo" nameprefix="" lastname="Magnini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:03:59.68">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2017-02-19" nation="ITA" />
     <ATHLETE firstname="Samuele" nameprefix="" lastname="Pampana" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:08:18.18">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Colle Val D&apos;Elsa" date="2016-02-06" nation="ITA" />
     <ATHLETE firstname="Samuele" nameprefix="" lastname="Pampana" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:15:51.60">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sori" date="2016-02-21" nation="ITA" />
     <ATHLETE firstname="Samuele" nameprefix="" lastname="Pampana" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:25.54">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Olsztyn" date="2018-11-17" nation="POL" />
     <ATHLETE firstname="Marcin" nameprefix="" lastname="Kaczmarek" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:00:56.22">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Padova" date="2023-03-19" nation="ITA" />
     <ATHLETE firstname="Enrico" nameprefix="" lastname="Catalano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:04.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Roma" date="2016-04-24" nation="ITA" />
     <ATHLETE firstname="Maurizio" nameprefix="" lastname="Tersar" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.68">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Funchal" date="2023-11-20" nation="POR" />
     <ATHLETE firstname="Filippo" nameprefix="" lastname="Magnini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:02.05">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2023-10-27" nation="GBR" />
     <ATHLETE firstname="Chris" nameprefix="" lastname="Jones" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:15.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Derby" date="2023-11-25" nation="GBR" />
     <ATHLETE firstname="Chris" nameprefix="" lastname="Jones" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:24.14">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sundsvall" date="2014-03-16" nation="SWE" />
     <ATHLETE firstname="Lars" nameprefix="" lastname="Fr�lander" gender="M" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:00:53.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sundsvall" date="2014-03-15" nation="SWE" />
     <ATHLETE firstname="Lars" nameprefix="" lastname="Fr�lander" gender="M" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:02:04.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Barcelona" date="2016-03-19" nation="ESP" />
     <ATHLETE firstname="Fernando" nameprefix="" lastname="Alaez" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:57.34">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2018-10-27" nation="GBR" />
     <ATHLETE firstname="Benjamin" nameprefix="" lastname="Harkin" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:06.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Troyes" date="2010-01-16" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:31.92">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Wuppertal" date="2011-11-05" nation="GER" />
     <ATHLETE firstname="Uwe" nameprefix="" lastname="Volk" gender="M" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:22.54">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-02-18" nation="" />
     <ATHLETE firstname="Mikel" nameprefix="" lastname="Bildosola Agirregomezkorta" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:49.64">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-06-04" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Hara" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:50.08">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2008-12-06" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Ross" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:00.67">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Bremen" date="2004-11-07" nation="GER" />
     <ATHLETE firstname="Kai" nameprefix="" lastname="Ditzel" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:08:15.69">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-02-25" nation="" />
     <ATHLETE firstname="Samuele" nameprefix="" lastname="Pampana" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:15:51.60">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-02-21" nation="" />
     <ATHLETE firstname="Samuele" nameprefix="" lastname="Pampana" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:25.48">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-03-21" nation="" />
     <ATHLETE firstname="M." nameprefix="" lastname="Wakabayashi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:54.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2008-12-07" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Ross" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:03.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2008-12-14" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Ross" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.06">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-12-05" nation="" />
     <ATHLETE firstname="Ryosuke" nameprefix="" lastname="Imai" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:01.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2014-12-06" nation="" />
     <ATHLETE firstname="Steven" nameprefix="" lastname="West" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:09.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-10-08" nation="" />
     <ATHLETE firstname="Brandon" nameprefix="" lastname="Fisher" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:23.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-10-01" nation="" />
     <ATHLETE firstname="Kohei" nameprefix="" lastname="Kawamoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:53.56">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-10-01" nation="" />
     <ATHLETE firstname="Kohei" nameprefix="" lastname="Kawamoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:02.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="1998-10-11" nation="" />
     <ATHLETE firstname="William" nameprefix="" lastname="Specht" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:56.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-03-19" nation="" />
     <ATHLETE firstname="Daisuke" nameprefix="" lastname="Hosokawa" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:03.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-12-02" nation="" />
     <ATHLETE firstname="Markus" nameprefix="" lastname="Rogan" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:30.68">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2014-10-10" nation="" />
     <ATHLETE firstname="Eric" nameprefix="" lastname="Christensen" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:24.22">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:00:52.71">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:02:01.79">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2009-11-29" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:27.04">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2008-02-02" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:09:25.61">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2007-01-20" nation="NED" />
     <ATHLETE firstname="Kees-Jan" nameprefix="van" lastname="Overbeeke" gender="M" nation="NED" CLUB="WWV Winterswijk" birthdate="1962-09-04" />
    </RECORD>
    <RECORD swimtime="00:18:13.37">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Winterswijk" date="2005-01-23" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:00:28.47">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Denekamp" date="2019-11-24" nation="NED" />
     <ATHLETE firstname="Tjakko" nameprefix="" lastname="Ruinemans" gender="M" nation="NED" CLUB="De Dinkel" birthdate="1974-08-23" />
    </RECORD>
    <RECORD swimtime="00:00:59.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Papendrecht" date="2009-11-29" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:12.87">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2008-03-16" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:30.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Arnhem" date="2013-03-16" nation="NED" />
     <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" CLUB="PSV" birthdate="1968-10-13" />
    </RECORD>
    <RECORD swimtime="00:01:08.83">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <ATHLETE firstname="Harry" nameprefix="" lastname="Cornet" gender="M" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1971-11-12" />
    </RECORD>
    <RECORD swimtime="00:02:29.71">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Vlijmen" date="2009-12-13" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:26.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:00:59.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:02:15.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Emmeloord" date="2006-01-21" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:00.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Papendrecht" date="2009-11-29" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:11.92">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Almere" date="2009-11-15" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:58.58">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2008-12-13" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:23.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Helsingborg" date="2016-05-07" nation="SWE" />
     <ATHLETE firstname="Joakim" nameprefix="" lastname="Holmquist" gender="M" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:00:51.30">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2012-03-10" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:52.87">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2012-03-09" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:03.10">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Trento" date="2015-04-18" nation="ITA" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:08:24.75">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rennes" date="2015-03-29" nation="FRA" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:16:08.41">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Livorno" date="2023-02-25" nation="ITA" />
     <ATHLETE firstname="Nicola" nameprefix="" lastname="Nisato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:25.73">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Poznan" date="2022-12-17" nation="POL" />
     <ATHLETE firstname="Marcin" nameprefix="" lastname="Kaczmarek" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:00:57.76">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Poznan" date="2022-12-17" nation="POL" />
     <ATHLETE firstname="Marcin" nameprefix="" lastname="Kaczmarek" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:02:06.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Angers" date="2012-03-11" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:28.87">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2010-01-17" nation="ITA" />
     <ATHLETE firstname="Rico" nameprefix="" lastname="Rolli" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:03.23">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rennes" date="2015-03-28" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:18.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rennes" date="2015-03-27" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:25.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Goslar" date="2023-03-04" nation="GER" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Herbst" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:56.37">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Angers" date="2016-03-25" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:07.50">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Mansea" date="2021-04-17" nation="ESP" />
     <ATHLETE firstname="Fernando" nameprefix="" lastname="Alaez" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:57.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Angers" date="2012-03-09" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:04.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Angers" date="2012-03-08" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:31.36">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Saint Dizier" date="2012-04-07" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:22.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-02-06" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Hara" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:49.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-02-06" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Hara" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:52.58">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-06-25" nation="" />
     <ATHLETE firstname="Rodrigo" nameprefix="" lastname="Castro" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:04:03.10">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-04-18" nation="" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:08:24.75">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-03-29" nation="" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:16:08.41">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-02-25" nation="" />
     <ATHLETE firstname="Nicola" nameprefix="" lastname="Nisato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:25.73">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-12-17" nation="" />
     <ATHLETE firstname="Marcin" nameprefix="" lastname="Kaczmarek" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:00:57.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2009-12-13" nation="" />
     <ATHLETE firstname="Chris" nameprefix="" lastname="Stevenson" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:05.54">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2009-12-12" nation="" />
     <ATHLETE firstname="Chris" nameprefix="" lastname="Stevenson" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.65">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-10-26" nation="" />
     <ATHLETE firstname="Jeff" nameprefix="" lastname="Commings" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:02.22">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-11-17" nation="" />
     <ATHLETE firstname="Steven" nameprefix="" lastname="West" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:15.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-11-30" nation="" />
     <ATHLETE firstname="Steven" nameprefix="" lastname="West" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:24.38">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-03-19" nation="" />
     <ATHLETE firstname="Eiji" nameprefix="" lastname="Nomura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:55.07">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2018-03-18" nation="" />
     <ATHLETE firstname="Eiji" nameprefix="" lastname="Nomura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:05.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2020-01-19" nation="" />
     <ATHLETE firstname="Eiji" nameprefix="" lastname="Nomura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:57.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Angers" date="2012-03-09" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:04.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Angers" date="2012-03-08" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:31.36">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2012-04-07" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:25.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-24" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:00:55.64">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1969-11-26" />
    </RECORD>
    <RECORD swimtime="00:02:04.85">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Nijverdal" date="2013-01-25" nation="NED" />
     <ATHLETE firstname="Cees" nameprefix="van" lastname="Houwelingen" gender="M" nation="NED" CLUB="De Schelde" birthdate="1963-03-24" />
    </RECORD>
    <RECORD swimtime="00:04:32.59">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-25" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:09:27.56">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <ATHLETE firstname="Bob" nameprefix="de" lastname="Vries" gender="M" nation="NED" CLUB="Aquapoldro" birthdate="1966-04-13" />
    </RECORD>
    <RECORD swimtime="00:18:10.09">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-19" nation="NED" />
     <ATHLETE firstname="Bob" nameprefix="de" lastname="Vries" gender="M" nation="NED" CLUB="Aquapoldro" birthdate="1966-04-13" />
    </RECORD>
    <RECORD swimtime="00:00:29.43">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1969-11-26" />
    </RECORD>
    <RECORD swimtime="00:01:01.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2014-06-28" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:16.23">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Zwolle" date="2014-01-26" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:31.63">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Arnhem" date="2018-03-24" nation="NED" />
     <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" CLUB="PSV" birthdate="1968-10-13" />
    </RECORD>
    <RECORD swimtime="00:01:10.61">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Arnhem" date="2018-03-24" nation="NED" />
     <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" CLUB="PSV" birthdate="1968-10-13" />
    </RECORD>
    <RECORD swimtime="00:02:33.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:26.97">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Vlissingen" date="2009-01-25" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:00:59.91">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Winterswijk" date="2008-05-03" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:12.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Vlaardingen" date="2010-01-22" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:01.21">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2014-07-05" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:17.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2015-01-23" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:58.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Vlissingen" date="2009-01-24" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:23.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eskilstuna" date="2019-03-23" nation="SWE" />
     <ATHLETE firstname="Joakim" nameprefix="" lastname="Holmquist" gender="M" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:00:51.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Dunkerque" date="2017-03-26" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:54.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Napoli" date="2018-05-05" nation="ITA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:04.48">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Cholet" date="2017-01-29" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:08:33.74">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vicenza" date="2018-11-17" nation="ITA" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:16:23.36">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Genova" date="2020-02-22" nation="ITA" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.13">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Gau-Algesheim" date="2023-01-14" nation="GER" />
     <ATHLETE firstname="Lars" nameprefix="" lastname="Kalenka" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:57.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Dunkerque" date="2017-03-25" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:07.13">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Giugliano" date="2017-05-06" nation="ITA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:29.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Istanbul" date="2023-08-26" nation="TUR" />
     <ATHLETE firstname="Serkan" nameprefix="" lastname="Atasay" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:01:04.28">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Giugliano" date="2017-05-06" nation="ITA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:19.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Angers" date="2018-03-23" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:25.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Mol" date="2023-03-25" nation="BEL" />
     <ATHLETE firstname="Fr�d�ric" nameprefix="" lastname="Tonus" gender="M" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:00:56.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Angers" date="2018-03-24" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:09.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Angers" date="2018-03-25" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:57.63">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Istanbul" date="2023-08-25" nation="TUR" />
     <ATHLETE firstname="Serkan" nameprefix="" lastname="Atasay" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:02:06.38">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Tours" date="2018-01-28" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:29.33">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Dunkerque" date="2017-03-23" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:23.36">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-05-28" nation="" />
     <ATHLETE firstname="Chris" nameprefix="" lastname="Fydler" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:00:51.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-03-26" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:54.61">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-10-14" nation="" />
     <ATHLETE firstname="Ambrose" nameprefix="" lastname="Gaines" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:04.48">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-01-29" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:08:33.74">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-11-17" nation="" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:16:23.36">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2020-02-22" nation="" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:26.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2015-10-24" nation="" />
     <ATHLETE firstname="Fritz" nameprefix="" lastname="Bedford" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:57.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-03-25" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:07.13">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-05-06" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:29.09">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-02-12" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Togo" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:04.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-02-12" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Togo" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:19.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-03-23" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:24.96">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-11-27" nation="JPN" />
     <ATHLETE firstname="Eiji" nameprefix="" lastname="Nomura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:55.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-01-15" nation="" />
     <ATHLETE firstname="Eiji" nameprefix="" lastname="Nomura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:07.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-01-15" nation="JPN" />
     <ATHLETE firstname="Eiji" nameprefix="" lastname="Nomura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:57.69">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-03-24" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:06.38">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-01-28" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:29.33">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-03-23" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:25.73">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:00:57.52">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2012-03-08" nation="FRA" />
     <ATHLETE firstname="Albert" nameprefix="" lastname="Boonstra" gender="M" nation="NED" CLUB="Aqua-Novio&apos;94" birthdate="1957-05-22" />
    </RECORD>
    <RECORD swimtime="00:02:05.07">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-24" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:04:30.73">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-25" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:09:23.27">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-26" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:18:12.52">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-24" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:00:29.49">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:01:03.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Terneuzen" date="2018-01-21" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:21.44">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Terneuzen" date="2018-01-21" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:32.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" CLUB="PSV" birthdate="1968-10-13" />
    </RECORD>
    <RECORD swimtime="00:01:12.67">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amsterdam" date="2008-02-16" nation="NED" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:02:39.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:27.35">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Nijverdal" date="2013-01-25" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:00.58">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Nijverdal" date="2013-01-27" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:15.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Nijverdal" date="2013-01-26" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:04.34">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2007-01-19" nation="NED" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:02:23.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Paris" date="2007-05-24" nation="FRA" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:02:23.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2015-01-23" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="Albion" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:05:07.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Nijverdal" date="2013-01-26" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:24.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-28" nation="GBR" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Hodgson" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:55.06">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Puy-en-Velay" date="2023-04-01" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:00.06">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Puy-en-Velay" date="2023-04-23" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:19.83">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2023-04-23" nation="ITA" />
     <ATHLETE firstname="Dino" nameprefix="" lastname="Schorn" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:09:01.71">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Torino" date="2023-02-12" nation="ITA" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:17:07.13">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Torino" date="2023-02-12" nation="ITA" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.96">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2016-10-30" nation="GBR" />
     <ATHLETE firstname="Craig" nameprefix="" lastname="Norrey" gender="M" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:01:02.26">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Trento" date="2015-03-15" nation="ITA" />
     <ATHLETE firstname="Marco" nameprefix="" lastname="Colombo" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:14.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Roma" date="2023-04-22" nation="ITA" />
     <ATHLETE firstname="Alessio" nameprefix="" lastname="Germani" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:29.22">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Lodi" date="2020-02-09" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:04.26">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Torino" date="2019-02-16" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:22.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2018-04-21" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:26.41">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Hannover" date="2023-12-02" nation="GER" />
     <ATHLETE firstname="Lars" nameprefix="" lastname="Renner" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:59.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Hannover" date="2023-12-02" nation="GER" />
     <ATHLETE firstname="Lars" nameprefix="" lastname="Renner" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:15.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Nijverdal" date="2013-01-26" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:01.28">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Guildford" date="2023-06-24" nation="GBR" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Hodgson" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:14.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Puy-en-Velay" date="2023-04-23" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:58.95">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Milano" date="2018-01-07" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:24.37">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-03-23" nation="" />
     <ATHLETE firstname="Calvin" nameprefix="" lastname="Maughan" gender="M" nation="rsa" />
    </RECORD>
    <RECORD swimtime="00:00:54.32">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-03-23" nation="" />
     <ATHLETE firstname="Calvin" nameprefix="" lastname="Maughan" gender="M" nation="rsa" />
    </RECORD>
    <RECORD swimtime="00:01:59.08">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-11-21" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:16.03">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-11-22" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:51.34">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-11-21" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:16:59.70">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-06-04" nation="" />
     <ATHLETE firstname="Brent" nameprefix="" lastname="Foster" gender="M" nation="NZL" />
    </RECORD>
    <RECORD swimtime="00:00:27.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-12-09" nation="" />
     <ATHLETE firstname="Fritz" nameprefix="" lastname="Bedford" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:00.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-10-20" nation="" />
     <ATHLETE firstname="Fritz" nameprefix="" lastname="Bedford" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:14.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-04-22" nation="" />
     <ATHLETE firstname="Alessio" nameprefix="" lastname="Germani" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:29.22">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2020-02-09" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:04.26">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-02-16" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:22.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-04-21" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:26.43">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-12-12" nation="" />
     <ATHLETE firstname="Steve" nameprefix="" lastname="Hiltabiddle" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:59.11">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-09-09" nation="" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Weldon" gender="M" nation="NZL" />
    </RECORD>
    <RECORD swimtime="00:02:15.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Nijverdal" date="2013-01-26" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:00.75">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-10-28" nation="" />
     <ATHLETE firstname="Mike" nameprefix="" lastname="Irvin" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:14.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-04-23" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:49.86">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-07-16" nation="" />
     <ATHLETE firstname="Brent" nameprefix="" lastname="Foster" gender="M" nation="NZL" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:26.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:00:59.27">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:02:11.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:04:40.45">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:09:44.41">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:18:47.47">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-18" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:00:30.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:08.48">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:02:29.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Vlaardingen" date="2022-12-11" nation="NED" />
     <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1962-02-13" />
    </RECORD>
    <RECORD swimtime="00:00:34.51">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2018-01-06" nation="NED" />
     <ATHLETE firstname="Albert" nameprefix="" lastname="Boonstra" gender="M" nation="NED" CLUB="Aqua-Novio&apos;94" birthdate="1957-05-22" />
    </RECORD>
    <RECORD swimtime="00:01:15.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amsterdam" date="2012-02-11" nation="NED" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:02:54.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2023-01-07" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:27.82">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="Feijenoord Albion zwemclub" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:01.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Terneuzen" date="2018-01-21" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:20.27">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:07.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Terneuzen" date="2012-01-28" nation="NED" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:02:26.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="Feijenoord Albion zwemclub" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:05:15.31">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Terneuzen" date="2018-01-21" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1958-09-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:25.37">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-21" nation="POR" />
     <ATHLETE firstname="Ahmet" nameprefix="" lastname="Nakkas" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:00:55.73">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-23" nation="POR" />
     <ATHLETE firstname="Ahmet" nameprefix="" lastname="Nakkas" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:02:05.16">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-20" nation="POR" />
     <ATHLETE firstname="Ahmet" nameprefix="" lastname="Nakkas" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:04:29.95">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Castellon" date="2023-02-17" nation="ESP" />
     <ATHLETE firstname="Juan Carlos" nameprefix="" lastname="Vallejo Arroyo" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:09:27.94">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Br�hl" date="2022-10-16" nation="GER" />
     <ATHLETE firstname="Karsten" nameprefix="" lastname="Dellbr�gge" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:18:23.61">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gau-Algesheim" date="2023-01-14" nation="GER" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Kleiber" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:29.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Plan-les-Oates" date="2022-03-31" nation="SUI" />
     <ATHLETE firstname="Craig" nameprefix="" lastname="Norrey" gender="M" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:01:05.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Poznan" date="2022-12-17" nation="POL" />
     <ATHLETE firstname="Zbigniew" nameprefix="" lastname="Korzeniowski" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:02:23.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Poznan" date="2022-12-18" nation="POL" />
     <ATHLETE firstname="Zbiegniew" nameprefix="" lastname="Korzeniowski" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:00:29.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2023-04-22" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:06.05">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Torino" date="2023-02-11" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:26.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2023-04-23" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="2022-10-30" nation="GBR" />
     <ATHLETE firstname="David" nameprefix="" lastname="Emerson" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:01.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Terneuzen" date="2018-01-21" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:20.27">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:03.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Lodi" date="2023-04-02" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:19.31">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Livorno" date="2023-02-25" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:05:05.11">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Paterno" date="2023-03-04" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:24.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2006-12-03" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:55.87">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-05-17" nation="" />
     <ATHLETE firstname="Jack" nameprefix="" lastname="Groselle" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:01.65">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-11-21" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:27.57">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-10-15" nation="" />
     <ATHLETE firstname="Arnaldo" nameprefix="" lastname="Perez" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:07.78">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-10-14" nation="" />
     <ATHLETE firstname="Arnaldo" nameprefix="" lastname="Perez" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:34.51">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-01-29" nation="" />
     <ATHLETE firstname="Arnaldo" nameprefix="" lastname="Perez" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:29.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-07-12" nation="" />
     <ATHLETE firstname="Jamie" nameprefix="" lastname="Fowler" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:03.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-07-12" nation="" />
     <ATHLETE firstname="Jamie" nameprefix="" lastname="Fowler" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:17.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-08-12" nation="" />
     <ATHLETE firstname="Jamie" nameprefix="" lastname="Fowler" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:29.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-04-22" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:06.05">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-02-11" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:26.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-04-23" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:26.78">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-05-13" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Thompson" gender="M" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:00.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2016-05-23" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Thompson" gender="M" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:02:20.27">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:03.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-04-02" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:19.31">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-02-25" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:05:04.54">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2011-11-13" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:27.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:01:00.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:16.33">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:04:50.72">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:09:58.48">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:19:29.25">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gouda" date="2023-03-12" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:00:33.54">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:10.02">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:35.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:00:36.51">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amsterdam" date="2019-05-25" nation="NED" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:01:19.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Papendrecht" date="2023-10-08" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:03:06.88">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2013-01-12" nation="NED" />
     <ATHLETE firstname="Donald" nameprefix="" lastname="Uijtenbogaart" gender="M" nation="NED" CLUB="Het Y" birthdate="1947-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:28.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:03.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:22.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:17.57">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2024-01-06" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:02:32.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:05:27.66">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2023-11-26" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:26.67">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Helsingb�rg" date="2016-05-07" nation="SWE" />
     <ATHLETE firstname="Leonard" nameprefix="" lastname="Bielicz" gender="M" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:01:00.37">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Helsingborg" date="2016-05-08" nation="SWE" />
     <ATHLETE firstname="Leonard" nameprefix="" lastname="Bielicz" gender="M" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:02:16.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2016-03-26" nation="FRA" />
     <ATHLETE firstname="Jean" nameprefix="Claude" lastname="Chatard" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:48.96">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2022-03-12" nation="FRA" />
     <ATHLETE firstname="Serge" nameprefix="" lastname="Guerin" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:09:58.48">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:19:21.87">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2018-03-24" nation="FRA" />
     <ATHLETE firstname="Patrick" nameprefix="" lastname="Moreau" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:31.91">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Boulogne" date="2019-04-06" nation="FRA" />
     <ATHLETE firstname="Pierre" nameprefix="" lastname="Baehr" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:09.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Angers" date="2022-03-10" nation="FRA" />
     <ATHLETE firstname="Jean" nameprefix="" lastname="Delaporte" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:35.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:33.88">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Palma de Mallorca" date="2019-04-27" nation="ESP" />
     <ATHLETE firstname="Pere" nameprefix="" lastname="Balcells Prat" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:16.34">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rennes" date="2015-03-28" nation="FRA" />
     <ATHLETE firstname="Christophe" nameprefix="" lastname="Starzec" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:50.38">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Birkesod" date="2021-03-13" nation="DEN" />
     <ATHLETE firstname="Sigitas" nameprefix="" lastname="Katkevicius" gender="M" nation="LTU" />
    </RECORD>
    <RECORD swimtime="00:00:28.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:03.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:22.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:08.72">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Papendrect" date="2023-10-08" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:32.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:05:27.66">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2023-11-26" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:25.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-03-03" nation="" />
     <ATHLETE firstname="Doug" nameprefix="" lastname="Martin" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:57.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-05-26" nation="" />
     <ATHLETE firstname="Jack" nameprefix="" lastname="Groselle" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:07.46">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-10-02" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Stephenson" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:27.91">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-11-19" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:26.94">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-11-24" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:18:26.04">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-06-23" nation="" />
     <ATHLETE firstname="Djan" nameprefix="" lastname="Garrido Madruga" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:00:30.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2012-12-02" nation="" />
     <ATHLETE firstname="Hugh" nameprefix="" lastname="Wilder" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:07.09">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-11-12" nation="" />
     <ATHLETE firstname="Jonathan" nameprefix="" lastname="Klein" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:28.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-04-02" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Stephenson" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:32.50">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-11-20" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:11.82">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-11-24" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:36.85">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-11-19" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:27.94">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-05-06" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Thompson" gender="M" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:03.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:22.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:01:05.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-11-19" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:20.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-11-17" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:03.34">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-11-18" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:30.41">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Reinier" nameprefix="" lastname="Dobbelmann" gender="M" nation="NED" CLUB="PSV" birthdate="1948-12-04" />
    </RECORD>
    <RECORD swimtime="00:01:09.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:02:33.73">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-10-31" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:05:30.15">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Grootebroek" date="2009-05-17" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:11:52.49">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vlissingen" date="2009-01-23" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:23:05.17">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vlaardingen" date="2010-01-22" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="De Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:00:35.71">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Hildesheim" date="2011-09-23" nation="GER" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:01:19.92">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:02:57.05">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:00:38.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Charles" nameprefix="" lastname="Bos" gender="M" nation="NED" CLUB="Patrick-De Roersoppers (SG)" birthdate="1953-05-22" />
    </RECORD>
    <RECORD swimtime="00:01:29.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Charles" nameprefix="" lastname="Bos" gender="M" nation="NED" CLUB="Patrick-De Roersoppers (SG)" birthdate="1953-05-22" />
    </RECORD>
    <RECORD swimtime="00:03:14.92">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Charles" nameprefix="" lastname="Bos" gender="M" nation="NED" CLUB="Patrick-De Roersoppers (SG)" birthdate="1953-05-22" />
    </RECORD>
    <RECORD swimtime="00:00:34.61">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:01:31.35">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Piet" nameprefix="" lastname="Schop" gender="M" nation="NED" CLUB="De Bevelanders" birthdate="1950-10-13" />
    </RECORD>
    <RECORD swimtime="00:03:33.94">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2008-03-16" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:01:22.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Charles" nameprefix="" lastname="Bos" gender="M" nation="NED" CLUB="Patrick-De Roersoppers (SG)" birthdate="1953-05-22" />
    </RECORD>
    <RECORD swimtime="00:03:15.01">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Almere-Stad" date="2008-11-23" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:07:02.20">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2013-02-16" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:28.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Link�ping" date="2008-03-08" nation="SWE" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bergengren" gender="M" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:01:03.91">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-23" nation="POR" />
     <ATHLETE firstname="Abed" nameprefix="" lastname="Ouadah" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:24.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-20" nation="POR" />
     <ATHLETE firstname="Abed" nameprefix="" lastname="Ouadah" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:05:07.58">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2022-03-12" nation="FRA" />
     <ATHLETE firstname="Patrick" nameprefix="" lastname="Moreau" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:10:32.27">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Angers" date="2022-03-10" nation="FRA" />
     <ATHLETE firstname="Patrick" nameprefix="" lastname="Moreau" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:20:45.27">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Glasgow" date="2023-11-04" nation="SCO" />
     <ATHLETE firstname="Eddie" nameprefix="" lastname="Riach" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:33.53">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Palma de Mallorca" date="2016-04-02" nation="ESP" />
     <ATHLETE firstname="Jean" nameprefix="" lastname="Lestideau" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:13.32">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Palma de Mallorca" date="2016-04-02" nation="ESP" />
     <ATHLETE firstname="Jean" nameprefix="" lastname="Lestideau" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:41.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Funchal" date="2023-11-23" nation="POR" />
     <ATHLETE firstname="Steve" nameprefix="" lastname="Grossman" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:35.53">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Villingen" date="2016-04-16" nation="GER" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="H�fer" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:22.45">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Villingen" date="2015-09-26" nation="GER" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="H�fer" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:05.27">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Gau Algesheim" date="2007-01-20" nation="GER" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Reichelt" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:31.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Oulu" date="2018-01-27" nation="FIN" />
     <ATHLETE firstname="Hannu" nameprefix="" lastname="Kuokkanen" gender="M" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:01:12.02">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2014-01-24" nation="NED" />
     <ATHLETE firstname="Josep" nameprefix="" lastname="Claret" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:53.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Dunkerque" date="2017-03-26" nation="FRA" />
     <ATHLETE firstname="Jean" nameprefix="" lastname="Lestideau" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:15.64">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Douglas" date="2018-02-17" nation="IRL" />
     <ATHLETE firstname="Kieran" nameprefix="" lastname="Kelleher" gender="M" nation="IRL" />
    </RECORD>
    <RECORD swimtime="00:02:43.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Angers" date="2022-03-13" nation="FRA" />
     <ATHLETE firstname="Patrick" nameprefix="" lastname="Moreau" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:05:46.48">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Angers" date="2022-03-10" nation="FRA" />
     <ATHLETE firstname="Patrick" nameprefix="" lastname="Moreau" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:26.88">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-10-10" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:01.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-05-17" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:01.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-01-22" nation="" />
     <ATHLETE firstname="Bruce" nameprefix="" lastname="Williams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:10.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-12-04" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:46.78">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-01-30" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:36.64">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-01-30" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:18:29.71">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-01-30" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:32.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-01-21" nation="USA" />
     <ATHLETE firstname="Bruce" nameprefix="" lastname="Williams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:11.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-11-13" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Day" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:34.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-11-14" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Day" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:33.54">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-12-04" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:13.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-12-04" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:55.87">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-03-05" nation="" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Strand" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:29.52">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2015-10-11" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:06.54">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-10-17" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Day" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:45.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-11-14" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Day" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:06.98">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-12-04" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:27.07">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-12-04" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:46.48">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-03-10" nation="" />
     <ATHLETE firstname="Patrick" nameprefix="" lastname="Moreau" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:33.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2014-02-09" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Z&amp;PC De Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:01:16.45">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2014-02-09" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Z&amp;PC De Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:02:51.74">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-24" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Z&amp;PC De Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:06:07.53">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2014-02-09" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Z&amp;PC De Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:13:13.28">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-18" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:24:53.01">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-18" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:00:37.87">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2015-01-24" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:01:24.58">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2015-01-24" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:03:03.13">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Heerenveen" date="2015-01-25" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:00:42.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Nijverdal" date="2013-01-26" nation="NED" />
     <ATHLETE firstname="Wieger" nameprefix="" lastname="Mensonides" gender="M" nation="NED" CLUB="NZ&amp;PC" birthdate="1938-07-12" />
    </RECORD>
    <RECORD swimtime="00:01:33.83">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Alphen a.d. Rijn" date="2018-02-18" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:03:28.89">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Paris" date="2018-08-05" nation="FRA" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:00:41.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2015-01-23" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:01:38.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Lelystad" date="2000-03-25" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:03:45.16">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Zwolle" date="2018-01-06" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:01:30.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Alphen a.d. Rijn" date="2018-02-18" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:03:22.04">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Alkmaar" date="2015-09-20" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:07:18.51">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Nijlen" date="2018-03-17" nation="BEL" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:29.47">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Graz" date="2019-02-09" nation="AUT" />
     <ATHLETE firstname="Gerhard" nameprefix="" lastname="Wieland" gender="M" nation="AUT" />
    </RECORD>
    <RECORD swimtime="00:01:07.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Hamburg-Dulsberg" date="2023-05-07" nation="GER" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="Seifert" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:34.44">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Hannover" date="2023-12-01" nation="GER" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="Seifert" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:05:44.36">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Palma de Mallorca" date="2016-04-02" nation="ESP" />
     <ATHLETE firstname="Joaquin " nameprefix="de" lastname="Canales Mendoza" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:12:03.35">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Bologna" date="2018-04-21" nation="ITA" />
     <ATHLETE firstname="Luciano" nameprefix="" lastname="Cammelli" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:23:18.51">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sabadell" date="2015-11-29" nation="ESP" />
     <ATHLETE firstname="Joaquin " nameprefix="de" lastname="Canales Mendoza" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:35.88">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Hamburg-Dulsberg" date="2023-05-07" nation="GER" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="Seifert" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:18.84">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Hamburg-Dulsberg" date="2023-05-07" nation="GER" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="Seifert" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:55.73">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Le Lamentin" date="2020-02-28" nation="FRA" />
     <ATHLETE firstname="Jozsef" nameprefix="" lastname="Csikany" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:00:36.78">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Lodi" date="2022-02-19" nation="ITA" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Rugieri" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:26.76">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Schweinfurt" date="2011-03-19" nation="GER" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Reichelt" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:15.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Schweinfurt" date="2011-03-20" nation="GER" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Reichelt" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:33.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sabadell" date="2020-01-12" nation="ESP" />
     <ATHLETE firstname="Josep" nameprefix="" lastname="Claret" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:19.34">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Goslar" date="2022-03-05" nation="GER" />
     <ATHLETE firstname="Horst" nameprefix="" lastname="Lehmann" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:10.85">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Ceska Lipa" date="2018-11-10" nation="CZE" />
     <ATHLETE firstname="Rudolf" nameprefix="" lastname="Smerda" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:20.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Hannover" date="2023-12-02" nation="GER" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="Seifert" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:00.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Hannover" date="2023-12-01" nation="GER" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="Seifert" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:06:33.07">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Allschwil" date="2021-10-31" nation="GER" />
     <ATHLETE firstname="Kurt" nameprefix="" lastname="Frei" gender="M" nation="SUI" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:28.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-11-21" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:04.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-10-13" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Quiggin" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:26.94">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-12-10" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Quiggin" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:09.95">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-03-11" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Kirkland" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:10:40.84">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-02-05" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Kirkland" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:20:18.58">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-02-05" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Kirkland" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:33.87">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-12-02" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:14.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-07-12" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:44.04">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-12-02" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:36.78">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-02-19" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Rugieri" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:24.27">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-12-03" nation="" />
     <ATHLETE firstname="Douglas" nameprefix="" lastname="Springer" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:06.82">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-07-23" nation="" />
     <ATHLETE firstname="Mike" nameprefix="" lastname="Freshley" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:32.09">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-11-21" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:17.51">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-10-29" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:10.85">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2018-11-10" nation="" />
     <ATHLETE firstname="Rudolf" nameprefix="" lastname="Smerda" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:17.58">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-07-23" nation="" />
     <ATHLETE firstname="Mike" nameprefix="" lastname="Freshley" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:50.79">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-11-30" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:26.09">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-09-22" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:36.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Winterswijk" date="2005-01-22" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:23.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2004-01-10" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:03:21.68">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vlaardingen" date="2022-12-11" nation="NED" />
     <ATHLETE firstname="G�za" nameprefix="" lastname="Kaltenecker" gender="M" nation="NED" CLUB="AZC" birthdate="1942-10-20" />
    </RECORD>
    <RECORD swimtime="00:07:04.19">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:14:57.64">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:29:18.23">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gouda" date="2023-03-12" nation="NED" />
     <ATHLETE firstname="G�za" nameprefix="" lastname="Kaltenecker" gender="M" nation="NED" CLUB="AZC" birthdate="1942-10-20" />
    </RECORD>
    <RECORD swimtime="00:00:43.54">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:01:32.98">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:03:33.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:00:45.82">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2004-01-10" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:50.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Winterswijk" date="2005-01-22" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:03:50.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2004-01-10" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:46.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Emmeloord" date="2006-01-22" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:43.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Heerenveen" date="2004-02-21" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:35.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2004-02-21" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:03:59.87">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Zwijndrecht" date="2023-04-08" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:09:26.59">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Barneveld" date="2024-01-20" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:32.07">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Wilhelmshaven" date="2019-01-26" nation="GER" />
     <ATHLETE firstname="Helmut" nameprefix="" lastname="Richter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:12.84">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Castellon" date="2012-01-27" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:45.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Castellon" date="2012-01-28" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:05:56.77">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Castellon" date="2012-01-28" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:12:50.20">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Fuengirola" date="2020-04-02" nation="ESP" />
     <ATHLETE firstname="Joaquin " nameprefix="de" lastname="Canales Mendoza" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:24:30.08">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Valladollid" date="2021-05-15" nation="ESP" />
     <ATHLETE firstname="Joaquin " nameprefix="de" lastname="Canales Mendoza" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:38.67">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Recklinghausen" date="2019-09-22" nation="GER" />
     <ATHLETE firstname="Helmut" nameprefix="" lastname="Richter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:21.74">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Funchal" date="2023-11-21" nation="POR" />
     <ATHLETE firstname="Jozsef" nameprefix="" lastname="Csikany" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:59.39">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Funchal" date="2023-11-23" nation="POR" />
     <ATHLETE firstname="Jozsef" nameprefix="" lastname="Csikany" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:00:42.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Innsbruck" date="2017-11-25" nation="AUT" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Reichelt" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:36.91">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Br�hl" date="2005-01-30" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:37.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Wilhelmshaven" date="2020-02-08" nation="GER" />
     <ATHLETE firstname="Joachim" nameprefix="" lastname="Schulze" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:35.98">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Palma de Mallorca" date="2024-01-20" nation="ESP" />
     <ATHLETE firstname="Josep" nameprefix="" lastname="Claret" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:30.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Genova" date="2011-12-03" nation="ITA" />
     <ATHLETE firstname="Giulio" nameprefix="" lastname="Divano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:03:30.11">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Genova" date="2011-02-27" nation="ITA" />
     <ATHLETE firstname="Giulio" nameprefix="" lastname="Divano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:28.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gau Algesheim" date="2015-01-18" nation="GER" />
     <ATHLETE firstname="Gerhard" nameprefix="" lastname="Hole" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:21.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Cadiz" date="2020-02-02" nation="ESP" />
     <ATHLETE firstname="Joaquin " nameprefix="de" lastname="Canales Mendoza" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:07:26.06">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Br�hl" date="2005-10-09" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:31.25">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-12-02" nation="" />
     <ATHLETE firstname="Jeff" nameprefix="" lastname="Farrell" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:09.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-02-12" nation="" />
     <ATHLETE firstname="Akira" nameprefix="" lastname="Fujimaki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:38.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-09-28" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:39.27">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-03-09" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:11:35.71">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-11-15" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:21:59.53">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-09-26" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:36.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-02-26" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:20.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-02-26" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:56.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-02-25" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:41.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2005-05-15" nation="" />
     <ATHLETE firstname="Toshio" nameprefix="" lastname="Tajima" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:31.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-02-21" nation="" />
     <ATHLETE firstname="Masaru" nameprefix="" lastname="Shinkai" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:21.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-02-21" nation="" />
     <ATHLETE firstname="Masaru" nameprefix="" lastname="Shinkai" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:34.92">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-02-25" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:29.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-09-02" nation="" />
     <ATHLETE firstname="Yasutaka" nameprefix="" lastname="Koike" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:30.11">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2011-02-27" nation="" />
     <ATHLETE firstname="Divano" nameprefix="" lastname="Giulio" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:23.73">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-02-26" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:08.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-02-25" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:07:09.74">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-04-15" nation="" />
     <ATHLETE firstname="Ikuro" nameprefix="" lastname="Shimono" gender="M" nation="JPN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:43.26">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gouda" date="2023-03-12" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:01:39.54">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gouda" date="2023-03-12" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:03:46.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:08:28.50">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" CLUB="PSV" birthdate="1933-04-17" />
    </RECORD>
    <RECORD swimtime="00:17:39.94">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-19" nation="POR" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:33:17.82">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gouda" date="2023-03-12" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:00:53.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="&apos;s-Gravenzande" date="2010-10-10" nation="NED" />
     <ATHLETE firstname="Ru" nameprefix="" lastname="Holtes" gender="M" nation="NED" CLUB="De Dolfijn" birthdate="1925-06-05" />
    </RECORD>
    <RECORD swimtime="00:01:59.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="&apos;s-Gravenzande" date="2010-10-10" nation="NED" />
     <ATHLETE firstname="Ru" nameprefix="" lastname="Holtes" gender="M" nation="NED" CLUB="De Dolfijn" birthdate="1925-06-05" />
    </RECORD>
    <RECORD swimtime="00:04:26.47">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Vlaardingen" date="2010-01-22" nation="NED" />
     <ATHLETE firstname="Ru" nameprefix="" lastname="Holtes" gender="M" nation="NED" CLUB="De Dolfijn" birthdate="1925-06-05" />
    </RECORD>
    <RECORD swimtime="00:01:13.17">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2013-01-12" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="00:02:59.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Zwolle" date="2014-01-26" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934 " birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:41.24">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" CLUB="PSV" birthdate="1933-04-17" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:32.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gijon" date="2016-01-29" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:14.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gijon" date="2016-01-31" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:55.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gijon" date="2016-01-30" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:06:30.16">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Malaga" date="2016-12-18" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:14:25.82">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <ATHLETE firstname="Frederik-Henrik" nameprefix="" lastname="De Bruijn" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:27:57.05">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Uimahalli" date="2022-03-25" nation="FIN" />
     <ATHLETE firstname="Lauri" nameprefix="" lastname="Malk" gender="M" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:00:43.83">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Gijon" date="2016-01-30" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:42.84">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Br�hl" date="2010-01-24" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:43.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Angers" date="2022-03-11" nation="FRA" />
     <ATHLETE firstname="Erwin" nameprefix="" lastname="Nodenschneider" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:45.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Innsbruck" date="2021-10-02" nation="AUT" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Reichelt" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:42.69">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Innsbruck" date="2021-10-03" nation="AUT" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Reichelt" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:55.71">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Manresa" date="2023-01-22" nation="ESP" />
     <ATHLETE firstname="Frederik-Henrik" nameprefix="" lastname="De Bruijn" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:41.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Gijon" date="2016-01-28" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:51.51">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Uimahalli" date="2022-03-27" nation="FIN" />
     <ATHLETE firstname="Lauri" nameprefix="" lastname="Malk" gender="M" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:04:07.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="2023-10-28" nation="GBR" />
     <ATHLETE firstname="David" nameprefix="" lastname="Cumming" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:34.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Murcia" date="2016-03-05" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:03:55.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Wuppertal" date="2011-11-05" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:08:08.28">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2023-10-27" nation="GBR" />
     <ATHLETE firstname="David" nameprefix="" lastname="Cumming" gender="M" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:32.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-01-29" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:14.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-01-31" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:55.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-01-30" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:06:27.44">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-04-13" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:13:20.46">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-01-13" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:25:18.19">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-12-04" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:40.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2009-04-19" nation="" />
     <ATHLETE firstname="Keijiro" nameprefix="" lastname="Nakamura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:28.98">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2008-05-18" nation="" />
     <ATHLETE firstname="Keijiro" nameprefix="" lastname="Nakamura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:18.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2008-04-20" nation="" />
     <ATHLETE firstname="Keijiro" nameprefix="" lastname="Nakamura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:44.47">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-06-13" nation="" />
     <ATHLETE firstname="Toshio" nameprefix="" lastname="Tajima" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:40.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-05-28" nation="" />
     <ATHLETE firstname="Tony" nameprefix="" lastname="Goodwin" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:03:44.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-04-22" nation="" />
     <ATHLETE firstname="Tony" nameprefix="" lastname="Goodwin" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:00:41.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2016-01-28" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:49.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-05-21" nation="" />
     <ATHLETE firstname="John" nameprefix="" lastname="Cocks" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:04:07.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-10-27" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Cumming" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:34.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Murcia" date="2016-03-05" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:03:36.41">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-05-22" nation="" />
     <ATHLETE firstname="John" nameprefix="" lastname="Cocks" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:07:58.08">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-05-20" nation="" />
     <ATHLETE firstname="John" nameprefix="" lastname="Cocks" gender="M" nation="AUS" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:01:28.89">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="00:03:23.03">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Emmeloord" date="2019-03-16" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="00:08:46.33">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Steenwijk" date="2021-09-30" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="00:18:26.92">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Steenwijk" date="2021-09-30" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:03.26">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Andel" date="2015-03-15" nation="NED" />
     <ATHLETE firstname="Ru" nameprefix="" lastname="Holtes" gender="M" nation="NED" CLUB="De Dolfijn" birthdate="1925-06-05" />
    </RECORD>
    <RECORD swimtime="00:02:29.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Grootebroek" date="2016-04-24" nation="NED" />
     <ATHLETE firstname="Ru" nameprefix="" lastname="Holtes" gender="M" nation="NED" CLUB="De Dolfijn" birthdate="1925-06-05" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:14.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Heerenveen" date="2019-02-16" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="00:05:17.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:00:43.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Br�hl" date="2015-01-25" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:35.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Br�hl" date="2015-10-11" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:27.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Hannover" date="2016-11-25" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:07:51.75">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Br�hl" date="2017-10-22" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:18:36.25">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Link�ping" date="2008-03-07" nation="SWE" />
     <ATHLETE firstname="Nils" nameprefix="" lastname="Ferm" gender="M" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:36:10.67">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2018-11-24" nation="GBr" />
     <ATHLETE firstname="Edward" nameprefix="" lastname="Hoy" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:53.24">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Deidesheim" date="2002-06-30" nation="GER" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Reinst�dler" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:58.74">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Freiburg" date="2015-11-29" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:20.68">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Wuppertal" date="2022-10-06" nation="GER" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Reinst�dler" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:51.68">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Br�hl" date="2015-10-11" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:56.64">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Gelsenkirchen" date="2015-11-07" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:21.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Giesing Harlaching" date="2016-11-12" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:54.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Essen" date="2021-11-27" nation="GER" />
     <ATHLETE firstname="Curt" nameprefix="" lastname="Zeiss" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:23.21">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Freiburg" date="2015-11-28" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="00:01:53.75">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Freiburg" date="2015-11-28" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:17.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Hannover" date="2016-11-25" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:00:40.93">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-02-07" nation="" />
     <ATHLETE firstname="Toshimi" nameprefix="" lastname="Inatomi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:35.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-10-11" nation="" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:27.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-11-25" nation="" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:07:42.61">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-10-23" nation="" />
     <ATHLETE firstname="Katsura" nameprefix="" lastname="Suzuki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:16:04.18">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-09-27" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:30:12.33">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-05-27" nation="" />
     <ATHLETE firstname="Katsura" nameprefix="" lastname="Suzuki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:52.40">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-05-14" nation="" />
     <ATHLETE firstname="Mampei" nameprefix="" lastname="Seino" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:47.66">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2006-05-14" nation="" />
     <ATHLETE firstname="Goro" nameprefix="" lastname="Kobayashi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:59.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2007-05-27" nation="" />
     <ATHLETE firstname="Goro" nameprefix="" lastname="Kobayashi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:49.58">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2015-06-07" nation="" />
     <ATHLETE firstname="Toshio" nameprefix="" lastname="Tajima" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:56.64">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2015-11-07" nation="" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:21.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-11-12" nation="" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:54.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-11-27" nation="" />
     <ATHLETE firstname="Curt" nameprefix="" lastname="Zeiss" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:16.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2018-06-10" nation="" />
     <ATHLETE firstname="G.da" nameprefix="" lastname="Silva" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:05:24.08">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2015-10-11" nation="" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Maine" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:53.75">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-11-28" nation="" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:17.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-11-25" nation="" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:09:39.56">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-11-15" nation="" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Maine" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:01:00.40">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gau Algesheim" date="2007-01-21" nation="GER" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Reinst�dler" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:36.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Castellon" date="2023-02-16" nation="ESP" />
     <ATHLETE firstname="Juan" nameprefix="" lastname="Dominguez" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:05:22.05">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Castellon" date="2023-02-18" nation="ESP" />
     <ATHLETE firstname="Juan" nameprefix="" lastname="Dominguez" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:10:39.55">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Pontevedra" date="2022-03-04" nation="ESP" />
     <ATHLETE firstname="Juan" nameprefix="" lastname="Dominguez" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:42:14.70">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Nyon" date="2019-11-02" nation="SUI" />
     <ATHLETE firstname="Werner" nameprefix="" lastname="Keller" gender="M" nation="SUI" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="00:01:03.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Gy�r" date="2015-04-12" nation="HUN" />
     <ATHLETE firstname="Bela Banki" nameprefix="" lastname="Horvath" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:29.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Gy�r" date="2015-04-11" nation="HUN" />
     <ATHLETE firstname="Bela Banki" nameprefix="" lastname="Horvath" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:06:18.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Isle of Wight" date="2009-02-22" nation="GBR" />
     <ATHLETE firstname="John" nameprefix="" lastname="Harrison" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:42.76">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Plan les Ouates" date="2019-04-06" nation="SUI" />
     <ATHLETE firstname="Werner" nameprefix="" lastname="Keller" gender="M" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:04:29.87">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Nyon" date="2019-12-08" nation="SUI" />
     <ATHLETE firstname="Werner" nameprefix="" lastname="Keller" gender="M" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:09:39.67">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Nyon" date="2019-11-02" nation="SUI" />
     <ATHLETE firstname="Werner" nameprefix="" lastname="Keller" gender="M" nation="SUI" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:00:45.47">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-11-18" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:47.23">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-03-04" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:56.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-11-18" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:13.42">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-03-05" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:16:56.22">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-11-19" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:31:56.67">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-11-19" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:55.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-11-19" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:04.72">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-11-11" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:24.83">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-11-18" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:07.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-01-24" nation="" />
     <ATHLETE firstname="Himoru" nameprefix="" lastname="Yoshimoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:31.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-01-24" nation="" />
     <ATHLETE firstname="Himoru" nameprefix="" lastname="Yoshimoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:05:45.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-05-08" nation="" />
     <ATHLETE firstname="Himoru" nameprefix="" lastname="Yoshimoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:02.24">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2018-10-27" nation="" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Doud" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:36.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2018-03-17" nation="" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Doud" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:11:08.68">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2018-03-17" nation="" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Doud" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:39.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-12-09" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:50.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2008-10-05" nation="" />
     <ATHLETE firstname="Walter" nameprefix="" lastname="Pfeiffer" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:21:03.17">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2008-10-05" nation="" />
     <ATHLETE firstname="Walter" nameprefix="" lastname="Pfeiffer" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="00:01:52.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Nogent sur Oise" date="2014-02-16" nation="FRA" />
     <ATHLETE firstname="Jean" nameprefix="" lastname="Leemput" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:03:33.45">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Godalming" date="2014-01-25" nation="GBR" />
     <ATHLETE firstname="John" nameprefix="" lastname="Harrison" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="00:01:26.68">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Paris" date="2014-03-29" nation="FRA" />
     <ATHLETE firstname="Jean" nameprefix="" lastname="Leemput" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:03:26.09">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Paris" date="2014-03-28" nation="FRA" />
     <ATHLETE firstname="Jean" nameprefix="" lastname="Leemput" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="00:00:55.75">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-06-23" nation="" />
     <ATHLETE firstname="George" nameprefix="" lastname="Corones" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:02:13.96">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-03-12" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:50.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-03-12" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:10:05.73">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-01-30" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:20:23.87">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-01-30" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:38:32.90">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-01-30" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:07.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-03-12" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:24.84">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-03-12" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:09.10">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-03-13" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:52.04">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-03-13" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="105" agemax="109" />
   <RECORDS>
    <RECORD swimtime="00:02:52.48">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-01-24" nation="" />
     <ATHLETE firstname="Jaring" nameprefix="" lastname="Timmerman" gender="M" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:03:09.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2014-01-24" nation="" />
     <ATHLETE firstname="Jaring" nameprefix="" lastname="Timmerman" gender="M" nation="CAN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="20" agemax="24" />
   <RECORDS>
    <RECORD swimtime="00:00:25.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="startlimiet" nameprefix="" lastname="" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:56.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Sam" nameprefix="van" lastname="Nunen" gender="F" nation="NED" CLUB="PSV" birthdate="2001-03-15" />
    </RECORD>
    <RECORD swimtime="00:02:07.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Sam" nameprefix="van" lastname="Nunen" gender="F" nation="NED" CLUB="PSV" birthdate="2001-03-15" />
    </RECORD>
    <RECORD swimtime="00:04:33.11">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-05-08" nation="NED" />
     <ATHLETE firstname="Marion" nameprefix="van den" lastname="Berg" gender="F" nation="NED" CLUB="DWK" birthdate="1986-01-01" />
    </RECORD>
    <RECORD swimtime="00:09:16.61">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-05-08" nation="NED" />
     <ATHLETE firstname="Marion" nameprefix="van den" lastname="Berg" gender="F" nation="NED" CLUB="DWK" birthdate="1986-01-01" />
    </RECORD>
    <RECORD swimtime="00:17:30.58">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-05-08" nation="NED" />
     <ATHLETE firstname="Marion" nameprefix="van den" lastname="Berg" gender="F" nation="NED" CLUB="DWK" birthdate="1986-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:29.64">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2014-05-03" nation="NED" />
     <ATHLETE firstname="Anja" nameprefix="van der" lastname="Hout" gender="F" nation="NED" CLUB="WVZ" birthdate="1990-06-18" />
    </RECORD>
    <RECORD swimtime="00:01:06.22">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Alkmaar" date="2018-04-08" nation="NED" />
     <ATHLETE firstname="Mirl" nameprefix="de" lastname="Boer" gender="F" nation="NED" CLUB="DAW" birthdate="1997-05-13" />
    </RECORD>
    <RECORD swimtime="00:02:24.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2012-05-04" nation="NED" />
     <ATHLETE firstname="Judith" nameprefix="van" lastname="Meijel" gender="F" nation="NED" CLUB="HZPC" birthdate="1991-06-26" />
    </RECORD>
    <RECORD swimtime="00:00:34.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="startlimiet" nameprefix="" lastname="" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:14.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Valesca" nameprefix="van den" lastname="Bogert" gender="F" nation="NED" CLUB="Hieronymus" birthdate="2001-04-06" />
    </RECORD>
    <RECORD swimtime="00:02:39.11">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Valesca" nameprefix="van den" lastname="Bogert" gender="F" nation="NED" CLUB="Hieronymus" birthdate="2001-04-06" />
    </RECORD>
    <RECORD swimtime="00:00:27.98">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Sam" nameprefix="van" lastname="Nunen" gender="F" nation="NED" CLUB="PSV" birthdate="2001-03-15" />
    </RECORD>
    <RECORD swimtime="00:01:03.54">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Luxembourg" date="2014-10-18" nation="LUX" />
     <ATHLETE firstname="Lisa" nameprefix="" lastname="Dreesens" gender="F" nation="NED" CLUB="PSV" birthdate="1991-10-05" />
    </RECORD>
    <RECORD swimtime="00:02:21.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="startlimiet" nameprefix="" lastname="" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:26.46">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2012-05-05" nation="NED" />
     <ATHLETE firstname="Wendan" nameprefix="" lastname="Poelstra" gender="F" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1991-09-15" />
    </RECORD>
    <RECORD swimtime="00:05:10.65">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Valesca" nameprefix="van den" lastname="Bogert" gender="F" nation="NED" CLUB="Hieronymus" birthdate="2001-04-06" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:25.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2004-02-15" nation="NED" />
     <ATHLETE firstname="Annabel" nameprefix="" lastname="Kosten" gender="F" nation="NED" CLUB="AZ&amp;PC" birthdate="1977-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:58.30">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Tamara" nameprefix="" lastname="Grove" gender="F" nation="NED" CLUB="De Dolfijn" birthdate="1996-10-02" />
    </RECORD>
    <RECORD swimtime="00:02:07.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Tamara" nameprefix="" lastname="Grove" gender="F" nation="NED" CLUB="De Dolfijn" birthdate="1996-10-02" />
    </RECORD>
    <RECORD swimtime="00:04:32.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Tamara" nameprefix="" lastname="Grove" gender="F" nation="NED" CLUB="De Dolfijn" birthdate="1996-10-02" />
    </RECORD>
    <RECORD swimtime="00:09:22.57">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Cadiz" date="2009-09-15" nation="ESP" />
     <ATHLETE firstname="Bianca" nameprefix="de" lastname="Bruijn" gender="F" nation="NED" CLUB="De Devel" birthdate="1984-11-09" />
    </RECORD>
    <RECORD swimtime="00:18:18.61">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-05" nation="NED" />
     <ATHLETE firstname="Lisa" nameprefix="" lastname="Dreesens" gender="F" nation="NED" CLUB="PSV" birthdate="1991-10-05" />
    </RECORD>
    <RECORD swimtime="00:00:30.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <ATHLETE firstname="Anja" nameprefix="van der" lastname="Hout" gender="F" nation="NED" CLUB="WVZ" birthdate="1990-06-18" />
    </RECORD>
    <RECORD swimtime="00:01:06.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <ATHLETE firstname="Anja" nameprefix="van der" lastname="Hout" gender="F" nation="NED" CLUB="WVZ" birthdate="1990-06-18" />
    </RECORD>
    <RECORD swimtime="00:02:23.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" CLUB="WVZ" birthdate="1993-11-05" />
    </RECORD>
    <RECORD swimtime="00:00:33.37">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-20" nation="HUN" />
     <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1988-07-28" />
    </RECORD>
    <RECORD swimtime="00:01:13.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2017-05-06" nation="NED" />
     <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1988-07-28" />
    </RECORD>
    <RECORD swimtime="00:02:44.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2017-05-05" nation="NED" />
     <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1988-07-28" />
    </RECORD>
    <RECORD swimtime="00:00:28.09">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Danique" nameprefix="" lastname="Stoop" gender="F" nation="NED" CLUB="Zuiderzeezwemmers" birthdate="1991-12-28" />
    </RECORD>
    <RECORD swimtime="00:01:03.01">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2017-03-26" nation="NED" />
     <ATHLETE firstname="Elinore" nameprefix="de" lastname="Jong" gender="F" nation="NED" CLUB="The Hague Swimming (SG)" birthdate="1989-04-23" />
    </RECORD>
    <RECORD swimtime="00:02:25.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Marlijn" nameprefix="" lastname="Hendriksen" gender="F" nation="NED" CLUB="Arethusa" birthdate="1988-08-16" />
    </RECORD>
    <RECORD swimtime="00:02:23.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Marjolein" nameprefix="" lastname="Delno" gender="F" nation="NED" CLUB="VZC" birthdate="1994-03-17" />
    </RECORD>
    <RECORD swimtime="00:05:18.38">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Budapest" date="2017-08-16" nation="HUN" />
     <ATHLETE firstname="Marlijn" nameprefix="" lastname="Hendriksen" gender="F" nation="NED" CLUB="Arethusa" birthdate="1988-08-16" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:25.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2004-02-15" nation="NED" />
     <ATHLETE firstname="Annabel" nameprefix="" lastname="Kosten" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:56.96">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kazan" date="2015-08-11" nation="RUS" />
     <ATHLETE firstname="Emma" nameprefix="" lastname="Gage" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:05.41">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2016-05-26" nation="GBR" />
     <ATHLETE firstname="Aisha" nameprefix="" lastname="Thornton" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:04:18.62">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Leeds" date="2011-06-18" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:45.89">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-12" nation="GER" />
     <ATHLETE firstname="Swann" nameprefix="" lastname="Oberson" gender="F" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:16:34.89">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-11" nation="GER" />
     <ATHLETE firstname="Swann" nameprefix="" lastname="Oberson" gender="F" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:00:29.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Roma" date="2022-08-30" nation="ITA" />
     <ATHLETE firstname="Valentina" nameprefix="" lastname="Catania" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:04.86">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Citavecchia" date="2021-07-03" nation="ITA" />
     <ATHLETE firstname="Valentina" nameprefix="" lastname="Catania" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:17.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Leeds" date="2011-06-18" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:32.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Pzmplona" date="1989-06-23" nation="ESP" />
     <ATHLETE firstname="Sabrina" nameprefix="" lastname="Seminatore" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:10.63">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="London" date="2016-05-27" nation="GBR" />
     <ATHLETE firstname="Rachael" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:35.82">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Cadiz" date="2009-09-19" nation="ESP" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:27.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Kazan" date="2015-08-12" nation="RUS" />
     <ATHLETE firstname="Emma" nameprefix="" lastname="Gage" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Kazan" date="2015-08-13" nation="RUS" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Polyakova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:18.77">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Mulhouse" date="2022-06-23" nation="FRA" />
     <ATHLETE firstname="Fanny" nameprefix="" lastname="Borer" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:21.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="St. Petersburg" date="2012-05-19" nation="RUS" />
     <ATHLETE firstname="Svetlana" nameprefix="" lastname="Karpeeva" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:05:04.80">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="K�ln" date="2015-04-18" nation="GER" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Spietzack" gender="F" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:25.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2004-02-15" nation="NED" />
     <ATHLETE firstname="Annabel" nameprefix="" lastname="Kosten" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:56.96">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-08-11" nation="" />
     <ATHLETE firstname="Emma" nameprefix="" lastname="Gage" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:04.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2010-07-10" nation="" />
     <ATHLETE firstname="Megan" nameprefix="" lastname="Jendrick" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:18.62">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Leeds" date="2011-06-18" nation="GBR" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:45.89">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2012-03-10" nation="" />
     <ATHLETE firstname="Swann" nameprefix="" lastname="Oberson" gender="F" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:16:34.89">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2012-03-11" nation="" />
     <ATHLETE firstname="Swann" nameprefix="" lastname="Oberson" gender="F" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:00:28.39">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-08-02" nation="" />
     <ATHLETE firstname="Emi" nameprefix="" lastname="Moronuki" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:01.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-07-31" nation="" />
     <ATHLETE firstname="Emi" nameprefix="" lastname="Moronuki" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:13.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-07-30" nation="" />
     <ATHLETE firstname="Emi" nameprefix="" lastname="Moronuki" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:31.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-07-10" nation="" />
     <ATHLETE firstname="Megan" nameprefix="" lastname="Jendrick" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:10.56">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-07-10" nation="" />
     <ATHLETE firstname="Megan" nameprefix="" lastname="Jendrick" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:32.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-06-24" nation="" />
     <ATHLETE firstname="Irina" nameprefix="" lastname="Shvaeva" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:26.32">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-06-16" nation="" />
     <ATHLETE firstname="Masako" nameprefix="" lastname="Kuroki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2015-08-13" nation="" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Polyakova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:15.02">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-05-20" nation="" />
     <ATHLETE firstname="Hannah" nameprefix="" lastname="Saiz" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:20.71">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2005-10-02" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:05:02.78">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2006-11-05" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:27.31">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <ATHLETE firstname="Pauline" nameprefix="" lastname="Gouwens" gender="F" nation="NED" CLUB="DWK" birthdate="1984-11-23" />
    </RECORD>
    <RECORD swimtime="00:00:59.16">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <ATHLETE firstname="Pauline" nameprefix="" lastname="Gouwens" gender="F" nation="NED" CLUB="DWK" birthdate="1984-11-23" />
    </RECORD>
    <RECORD swimtime="00:02:08.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" CLUB="WVZ" birthdate="1993-11-05" />
    </RECORD>
    <RECORD swimtime="00:04:36.20">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" CLUB="WVZ" birthdate="1993-11-05" />
    </RECORD>
    <RECORD swimtime="00:09:35.48">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" CLUB="WVZ" birthdate="1993-11-05" />
    </RECORD>
    <RECORD swimtime="00:18:48.96">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2012-05-04" nation="NED" />
     <ATHLETE firstname="Ann" nameprefix="" lastname="Wanter" gender="F" nation="NED" CLUB="Orca" birthdate="1982-10-29" />
    </RECORD>
    <RECORD swimtime="00:00:31.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <ATHLETE firstname="Evy" nameprefix="" lastname="Witlox" gender="F" nation="NED" CLUB="DWT" birthdate="1988-08-28" />
    </RECORD>
    <RECORD swimtime="00:01:08.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Evy" nameprefix="" lastname="Witlox" gender="F" nation="NED" CLUB="DWT" birthdate="1988-08-28" />
    </RECORD>
    <RECORD swimtime="00:02:23.47">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kiel" date="1993-04-24" nation="GER" />
     <ATHLETE firstname="Daphne" nameprefix="" lastname="Fuchs-Demuth" gender="F" nation="NED" CLUB="SG Minden-Porta" birthdate="1962-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:33.15">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1988-07-28" />
    </RECORD>
    <RECORD swimtime="00:01:13.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1988-07-28" />
    </RECORD>
    <RECORD swimtime="00:02:44.98">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Loes" nameprefix="" lastname="Zanderink" gender="F" nation="NED" CLUB="SwimGym" birthdate="1988-11-23" />
    </RECORD>
    <RECORD swimtime="00:00:28.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Danique" nameprefix="" lastname="Stoop" gender="F" nation="NED" CLUB="Zuiderzeezwemmers" birthdate="1991-12-28" />
    </RECORD>
    <RECORD swimtime="00:01:04.23">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <ATHLETE firstname="Elinore" nameprefix="de" lastname="Jong" gender="F" nation="NED" CLUB="The Hague Swimming (SG)" birthdate="1989-04-23" />
    </RECORD>
    <RECORD swimtime="00:02:29.65">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Marlijn" nameprefix="" lastname="Hendriksen" gender="F" nation="NED" CLUB="Hieronymus" birthdate="1988-08-16" />
    </RECORD>
    <RECORD swimtime="00:02:29.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Christchurch" date="2002-03-24" nation="NZL" />
     <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" CLUB="AZ&amp;PC" birthdate="1970-07-01" />
    </RECORD>
    <RECORD swimtime="00:05:17.89">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Marlijn" nameprefix="" lastname="Hendriksen" gender="F" nation="NED" CLUB="Hieronymus" birthdate="1988-08-16" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:26.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kazan" date="2015-08-14" nation="RUS" />
     <ATHLETE firstname="Irina" nameprefix="" lastname="Shlemova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:57.65">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kazan" date="2015-08-11" nation="RUS" />
     <ATHLETE firstname="Irina" nameprefix="" lastname="Shlemova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:05.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sydney" date="2013-04-18" nation="AUS" />
     <ATHLETE firstname="Caroline" nameprefix="" lastname="Saxby" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:04:22.91">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-20" nation="HUN" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:58.94">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-14" nation="HUN" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:17:20.55">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Aberdeen" date="2017-06-16" nation="SCO" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:29.49">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Aqua City" date="2023-09-24" nation="RUS" />
     <ATHLETE firstname="Anastasiya" nameprefix="" lastname="Fesikova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:03.30">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Crawley" date="2012-01-29" nation="GBR" />
     <ATHLETE firstname="Katy" nameprefix="" lastname="Sexton" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:18.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Aberdeen" date="2017-06-18" nation="SCO" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:31.88">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kranj" date="2018-09-03" nation="SLO" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Chocova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:11.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kazan" date="2015-08-11" nation="RUS" />
     <ATHLETE firstname="Natalia" nameprefix="" lastname="Vinokourenkova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:35.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Montreal" date="2014-08-08" nation="CAN" />
     <ATHLETE firstname="Natalia" nameprefix="" lastname="Vinokourenkova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:27.75">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Gwangju" date="2019-08-14" nation="KOR" />
     <ATHLETE firstname="Suvi" nameprefix="" lastname="Pulkkinen" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:01:01.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-08" nation="JPN" />
     <ATHLETE firstname="Afroditi" nameprefix="" lastname="Giareni" gender="F" nation="GRE" />
    </RECORD>
    <RECORD swimtime="00:02:18.21">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-10" nation="JPN" />
     <ATHLETE firstname="Afroditi" nameprefix="" lastname="Giareni" gender="F" nation="GRE" />
    </RECORD>
    <RECORD swimtime="00:02:20.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Fukuoka" date="2023-08-08" nation="JPN" />
     <ATHLETE firstname="Afroditi" nameprefix="" lastname="Giareni" gender="F" nation="GRE" />
    </RECORD>
    <RECORD swimtime="00:05:02.23">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Montreal" date="2014-08-05" nation="CAN" />
     <ATHLETE firstname="Natalia" nameprefix="" lastname="Vinokourenkova" gender="F" nation="RUS" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:25.74">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Austin" date="2008-06-06" nation="USA" />
     <ATHLETE firstname="Martina" nameprefix="" lastname="Moravcova" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:55.24">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-07-11" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Erndl" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:02.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-08-14" nation="" />
     <ATHLETE firstname="Natthanan" nameprefix="" lastname="Junkrajang" gender="F" nation="THA" />
    </RECORD>
    <RECORD swimtime="00:04:18.63">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-07-16" nation="" />
     <ATHLETE firstname="Dawn" nameprefix="" lastname="Heckman" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:46.47">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-07-14" nation="" />
     <ATHLETE firstname="Dawn" nameprefix="" lastname="Heckman" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:20.55">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-06-16" nation="" />
     <ATHLETE firstname="Sophie" nameprefix="" lastname="Casson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:28.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2012-08-07" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:01.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2011-08-06" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:17.61">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2009-08-06" nation="" />
     <ATHLETE firstname="Sarabeth" nameprefix="" lastname="Metzger" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:32.22">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-09-03" nation="NED" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:10.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2009-10-03" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:28.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2009-10-17" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:27.48">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2008-06-07" nation="" />
     <ATHLETE firstname="Martina" nameprefix="" lastname="Moravcova" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:58.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2008-06-07" nation="" />
     <ATHLETE firstname="Martina" nameprefix="" lastname="Moravcova" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:13.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2006-05-07" nation="" />
     <ATHLETE firstname="Mette" nameprefix="" lastname="Jacobsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:02:13.89">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-07-07" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Erndl" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:56.08">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-11-08" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:28.31">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2012-05-06" nation="NED" />
     <ATHLETE firstname="Janneke" nameprefix="" lastname="Harmsen-Bakker" gender="F" nation="NED" CLUB="De Spatters" birthdate="1977-06-26" />
    </RECORD>
    <RECORD swimtime="00:01:01.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kranj" date="2018-09-06" nation="SLO" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:15.03">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-16" nation="HUN" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:04:49.20">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2008-01-19" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Het Y" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:09:50.01">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2008-01-20" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Het Y" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:18:37.27">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2007-04-22" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Het Y" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:00:33.00">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2012-05-06" nation="NED" />
     <ATHLETE firstname="Janneke" nameprefix="" lastname="Harmsen-Bakker" gender="F" nation="NED" CLUB="De Spatters" birthdate="1977-06-26" />
    </RECORD>
    <RECORD swimtime="00:01:11.97">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Wachtebeke" date="2023-03-04" nation="BEL" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Schouten" gender="F" nation="NED" CLUB="MZ&amp;PC" birthdate="1987-09-08" />
    </RECORD>
    <RECORD swimtime="00:02:38.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Munchen" date="2000-08-01" nation="GER" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Cromjongh" gender="F" nation="NED" CLUB="De Zwoer" birthdate="1964-03-17" />
    </RECORD>
    <RECORD swimtime="00:00:35.24">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-20" nation="HUN" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="DAW" birthdate="1982-04-05" />
    </RECORD>
    <RECORD swimtime="00:01:18.61">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Dani�lle" nameprefix="" lastname="Reijnders" gender="F" nation="NED" CLUB="AquAmigos" birthdate="1985-07-20" />
    </RECORD>
    <RECORD swimtime="00:02:52.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="DAW" birthdate="1982-04-05" />
    </RECORD>
    <RECORD swimtime="00:00:29.75">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:01:08.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-17" nation="HUN" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:37.88">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Roos" nameprefix="van" lastname="Esch" gender="F" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1982-07-17" />
    </RECORD>
    <RECORD swimtime="00:02:33.98">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:05:39.61">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2014-05-04" nation="NED" />
     <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" CLUB="PSV" birthdate="1975-03-04" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:26.58">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2017-07-01" nation="ITA" />
     <ATHLETE firstname="Olessia" nameprefix="" lastname="Bourova" gender="F" nation="ita" />
    </RECORD>
    <RECORD swimtime="00:00:58.22">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Girona" date="2015-05-09" nation="ESP" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Roca" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:09.58">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2016-05-26" nation="GBR" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Roca" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:04:34.48">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2022-08-29" nation="ITA" />
     <ATHLETE firstname="Anna" nameprefix="" lastname="Spietzack" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:09:20.69">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="roma" date="2022-08-28" nation="ITA" />
     <ATHLETE firstname="Maren" nameprefix="" lastname="Spietzack" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:17:57.14">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2017-03-04" nation="GBR" />
     <ATHLETE firstname="Emma" nameprefix="" lastname="Wills" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:30.47">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Budapest" date="2017-08-20" nation="HUN" />
     <ATHLETE firstname="Alena" nameprefix="" lastname="Nyvltova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:07.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2023-06-02" nation="GBR" />
     <ATHLETE firstname="victoria" nameprefix="" lastname="Reading" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:23.47">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Glasgow" date="2005-06-03" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:31.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Fukuoka" date="2023-08-11" nation="JPN" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Weber" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:11.01">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Fukuoka" date="2023-08-06" nation="JPN" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Weber" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:38.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:28.03">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-07" nation="JPN" />
     <ATHLETE firstname="Petra" nameprefix="" lastname="Weber" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:05.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-17" nation="HUN" />
     <ATHLETE firstname="Gabriela" nameprefix="" lastname="Kostkova" gender="F" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:23.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2022-09-02" nation="ITA" />
     <ATHLETE firstname="Vikt�ria" nameprefix="" lastname="H�den-Felf�ldi" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:25.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Kranj" date="2018-09-05" nation="SLO" />
     <ATHLETE firstname="Natalia" nameprefix="" lastname="Vinokourenkova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:05:10.13">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Silingen" date="2022-03-19" nation="GER" />
     <ATHLETE firstname="Maren" nameprefix="" lastname="Spietzack" gender="F" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:25.98">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2006-08-08" nation="" />
     <ATHLETE firstname="Dara" nameprefix="" lastname="Torres" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:57.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-12-01" nation="" />
     <ATHLETE firstname="Veronica" nameprefix="" lastname="Balsano" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:02:05.50">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-12-02" nation="" />
     <ATHLETE firstname="Veronica" nameprefix="" lastname="Balsano" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:04:26.17">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="1997-08-10" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:09:08.47">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2012-11-18" nation="" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:17:17.22">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-08-06" nation="" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.63">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2016-08-18" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:01.75">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-08-19" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:18.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="1997-08-10" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:31.35">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-08-07" nation="" />
     <ATHLETE firstname="Danielle" nameprefix="" lastname="Herrmann" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:10.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-08-05" nation="" />
     <ATHLETE firstname="Danielle" nameprefix="" lastname="Herrmann" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:35.40">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2012-06-10" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:27.46">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2014-08-05" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:02.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-07-30" nation="" />
     <ATHLETE firstname="Carolina" nameprefix="" lastname="Sarruf" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:02:20.21">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="1997-08-10" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:21.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-08-06" nation="" />
     <ATHLETE firstname="Danielle" nameprefix="" lastname="Herrmann" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:59.59">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2012-06-16" nation="" />
     <ATHLETE firstname="Hitomi" nameprefix="" lastname="Matsuda" gender="F" nation="JPN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:26.64">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-09-06" nation="NED" />
     <ATHLETE firstname="Inge" nameprefix="de" lastname="Bruijn" gender="F" nation="NED" CLUB="PSV" birthdate="1973-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:01.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rome" date="2022-09-04" nation="ITA" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:02:17.92">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:04:49.48">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2012-05-05" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:09:52.17">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2012-05-06" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:18:47.76">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2012-05-04" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:00:33.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2012-05-05" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:01:13.56">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:02:40.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2013-09-05" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:00:35.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rome" date="2022-09-02" nation="ITA" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="DAW" birthdate="1982-04-05" />
    </RECORD>
    <RECORD swimtime="00:01:20.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="DAW" birthdate="1982-04-05" />
    </RECORD>
    <RECORD swimtime="00:02:53.58">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="DAW" birthdate="1982-04-05" />
    </RECORD>
    <RECORD swimtime="00:00:29.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Rome" date="2022-09-01" nation="ITA" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:01:08.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Cadiz" date="2009-09-16" nation="ESP" />
     <ATHLETE firstname="Anita" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="DIO" birthdate="1969-10-12" />
    </RECORD>
    <RECORD swimtime="00:02:37.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="G�teborg" date="2010-08-05" nation="SWE" />
     <ATHLETE firstname="Anita" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="DIO" birthdate="1969-10-12" />
    </RECORD>
    <RECORD swimtime="00:02:34.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" CLUB="WVZ" birthdate="1980-02-29" />
    </RECORD>
    <RECORD swimtime="00:05:38.89">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2010-05-07" nation="NED" />
     <ATHLETE firstname="Anita" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="DIO" birthdate="1969-10-12" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:26.64">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-09-06" nation="NED" />
     <ATHLETE firstname="Inge" nameprefix="de" lastname="Bruijn" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:59.63">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2016-05-28" nation="GBR" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:02:09.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-07" nation="NED" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:04:28.24">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Manchester" date="2015-06-14" nation="GBR" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:09:06.86">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Manchester" date="2015-06-12" nation="GBR" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:17:31.51">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2015-05-10" nation="NED" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:30.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="London" date="2016-05-27" nation="GBR" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:01:06.32">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:02:27.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Glasgow" date="2010-06-20" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:32.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2022-09-02" nation="ITA" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:12.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Berlin" date="2022-03-12" nation="GER" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:39.11">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2022-02-01" nation="ITA" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:28.68">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-16" nation="HUN" />
     <ATHLETE firstname="Raakel" nameprefix="" lastname="Luoto" gender="F" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:01:03.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Las Palmas" date="2022-07-11" nation="ESP" />
     <ATHLETE firstname="Mireia" nameprefix="" lastname="Garcia Sanchez" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:26.65">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Kinczo" nameprefix="" lastname="Venczel" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:26.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gwangju" date="2019-08-15" nation="KOR" />
     <ATHLETE firstname="Smiljana" nameprefix="" lastname="Marinovic" gender="F" nation="CRO" />
    </RECORD>
    <RECORD swimtime="00:05:15.53">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Valencia" date="2021-07-12" nation="ESP" />
     <ATHLETE firstname="Mirea" nameprefix="" lastname="Garcia" gender="F" nation="ESP" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:26.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-11-07" nation="" />
     <ATHLETE firstname="Edith" nameprefix="" lastname="Ottermann" gender="F" nation="RSA" />
    </RECORD>
    <RECORD swimtime="00:00:58.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-06-08" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:09.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2005-08-15" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:22.87">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-08-13" nation="" />
     <ATHLETE firstname="Janet" nameprefix="" lastname="Evans" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:59.06">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-06-11" nation="" />
     <ATHLETE firstname="Janet" nameprefix="" lastname="Evans" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:29.43">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-06-30" nation="" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:29.62">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-08-02" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:04.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-07-31" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:23.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2009-08-06" nation="" />
     <ATHLETE firstname="Jody" nameprefix="" lastname="Smith" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:32.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-09-02" nation="" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:12.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-03-12" nation="" />
     <ATHLETE firstname="Nicole" nameprefix="" lastname="Heidemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:38.44">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2006-08-09" nation="" />
     <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.36">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2013-06-08" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:03.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2009-05-23" nation="" />
     <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:24.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2006-07-23" nation="" />
     <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:25.03">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2007-08-05" nation="" />
     <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:09.83">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2004-08-01" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:28.00">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-04" nation="NED" />
     <ATHLETE firstname="Monique" nameprefix="" lastname="Tuijp" gender="F" nation="NED" CLUB="WZ&amp;PC Purmerend" birthdate="1969-01-28" />
    </RECORD>
    <RECORD swimtime="00:01:02.52">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" CLUB="PSV" birthdate="1973-11-06" />
    </RECORD>
    <RECORD swimtime="00:02:12.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" CLUB="PSV" birthdate="1973-11-06" />
    </RECORD>
    <RECORD swimtime="00:04:56.23">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" CLUB="PSV" birthdate="1975-03-04" />
    </RECORD>
    <RECORD swimtime="00:10:10.33">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-03" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="ZPCH" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:19:10.33">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-03" nation="NED" />
     <ATHLETE firstname="Grith" nameprefix="" lastname="Sigsgaard" gender="F" nation="NED" CLUB="ZPCH" birthdate="1972-09-25" />
    </RECORD>
    <RECORD swimtime="00:00:34.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:01:14.06">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:02:39.08">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1972-03-08" />
    </RECORD>
    <RECORD swimtime="00:00:36.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2017-05-07" nation="NED" />
     <ATHLETE firstname="Marjo" nameprefix="" lastname="Goelema-Koek" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1969-01-02" />
    </RECORD>
    <RECORD swimtime="00:01:21.14">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2017-05-06" nation="NED" />
     <ATHLETE firstname="Marjo" nameprefix="" lastname="Goelema-Koek" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1969-01-02" />
    </RECORD>
    <RECORD swimtime="00:02:59.16">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2007-04-20" nation="NED" />
     <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" CLUB="AZ&amp;PC" birthdate="1961-07-26" />
    </RECORD>
    <RECORD swimtime="00:00:30.94">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Aberdeen" date="2017-06-18" nation="GBR" />
     <ATHLETE firstname="Jeanne" nameprefix="" lastname="Petit" gender="F" nation="NED" CLUB="De Dinkel" birthdate="1970-02-13" />
    </RECORD>
    <RECORD swimtime="00:01:09.96">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2013-09-03" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="Neptunus" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:02:46.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2020-12-10" nation="NED" />
     <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" CLUB="PSV" birthdate="1975-03-04" />
    </RECORD>
    <RECORD swimtime="00:02:40.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1972-03-08" />
    </RECORD>
    <RECORD swimtime="00:05:43.75">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1972-03-08" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:27.04">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Antibes" date="2013-06-23" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:59.94">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="L�beck" date="2014-05-03" nation="GER" />
     <ATHLETE firstname="Barbara" nameprefix="" lastname="Kehbein" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:12.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:04:38.49">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2022-08-29" nation="ITA" />
     <ATHLETE firstname="Tiziana" nameprefix="" lastname="Papandrea" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:09:37.20">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Brescia" date="2016-03-05" nation="ITA" />
     <ATHLETE firstname="Valeria" nameprefix="" lastname="Vergani" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:18:33.06">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2023-03-04" nation="GBR" />
     <ATHLETE firstname="Ceri" nameprefix="" lastname="Edwards" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:31.58">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Budapest" date="2017-08-20" nation="HUN" />
     <ATHLETE firstname="Andrea" nameprefix="" lastname="Kutz" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:07.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Swansea" date="2019-06-14" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:24.06">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="London" date="2016-05-28" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:34.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Cadiz" date="2009-09-16" nation="ESP" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:13.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Cadiz" date="2009-09-17" nation="ESP" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:40.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Cadiz" date="2009-09-19" nation="ESP" />
     <ATHLETE firstname="Marzena" nameprefix="" lastname="Kulis" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:29.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Plymouth" date="2018-06-09" nation="GBR" />
     <ATHLETE firstname="Michelle" nameprefix="" lastname="Ware" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:06.91">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Riccione" date="2014-06-25" nation="ITA" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:27.71">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2019-04-14" nation="HUN" />
     <ATHLETE firstname="Kinczo" nameprefix="" lastname="Venczel" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:32.02">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="L�beck" date="2015-03-07" nation="GER" />
     <ATHLETE firstname="Barbara" nameprefix="" lastname="Kehbein" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:05:32.69">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="K�ln" date="2012-04-20" nation="GER" />
     <ATHLETE firstname="Angela" nameprefix="" lastname="Delissen" gender="F" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:26.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-03-16" nation="" />
     <ATHLETE firstname="Edith" nameprefix="" lastname="Ottermann" gender="F" nation="RSA" />
    </RECORD>
    <RECORD swimtime="00:00:57.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-08-08" nation="" />
     <ATHLETE firstname="Melanie" nameprefix="" lastname="Thomas" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:10.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-06-13" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:30.64">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-04-14" nation="" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:11.47">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-06-27" nation="" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:27.11">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-04-13" nation="" />
     <ATHLETE firstname="Heidi" nameprefix="" lastname="George" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:31.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2016-08-18" nation="" />
     <ATHLETE firstname="Cindy" nameprefix="" lastname="Mabee" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:07.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-06-14" nation="" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:24.06">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2016-05-28" nation="" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:33.56">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-08-20" nation="" />
     <ATHLETE firstname="Linley" nameprefix="" lastname="Frame" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:12.34">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-08-14" nation="" />
     <ATHLETE firstname="Gabrielle" nameprefix="" lastname="Rose" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:39.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-06-24" nation="" />
     <ATHLETE firstname="Gabrielle" nameprefix="" lastname="Rose" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.40">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-08-05" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:04.96">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2014-08-06" nation="" />
     <ATHLETE firstname="Wenke" nameprefix="" lastname="Seider" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:24.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2009-06-20" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:21.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-08-14" nation="" />
     <ATHLETE firstname="Gabrielle" nameprefix="" lastname="Rose" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:13.85">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2008-09-05" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:29.31">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:01:04.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg/Hollerich" date="2022-10-08" nation="LUX" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:02:20.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:04:52.14">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg/Hollerich" date="2022-10-08" nation="LUX" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:10:05.71">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:19:22.87">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-04" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:00:34.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:01:14.26">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:02:43.59">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" CLUB="PSV" birthdate="1972-02-07" />
    </RECORD>
    <RECORD swimtime="00:00:36.36">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kampen" date="2011-04-16" nation="NED" />
     <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" CLUB="AZ&amp;PC" birthdate="1961-07-26" />
    </RECORD>
    <RECORD swimtime="00:01:22.58">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-09-04" nation="NED" />
     <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" CLUB="AZ&amp;PC" birthdate="1961-07-26" />
    </RECORD>
    <RECORD swimtime="00:03:02.10">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kampen" date="2011-04-16" nation="NED" />
     <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" CLUB="AZ&amp;PC" birthdate="1961-07-26" />
    </RECORD>
    <RECORD swimtime="00:00:31.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:01:12.61">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2009-08-23" nation="NED" />
     <ATHLETE firstname="Mathilde" nameprefix="" lastname="Vink" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1958-12-12" />
    </RECORD>
    <RECORD swimtime="00:02:41.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:02:45.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
    <RECORD swimtime="00:05:38.55">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Luxembourg/Hollerich" date="2022-10-08" nation="LUX" />
     <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1971-04-20" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:27.09">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Chalon" date="2015-06-28" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:00.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Chalon" date="2015-06-27" nation="FRA" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:16.01">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Zaragoza" date="2015-07-24" nation="ESP" />
     <ATHLETE firstname="Maria" nameprefix="" lastname="Garcia" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:04:42.89">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Scanzano" date="2023-06-11" nation="ITA" />
     <ATHLETE firstname="Tiziana" nameprefix="" lastname="Papandrea" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:09:40.01">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2023-06-27" nation="ITA" />
     <ATHLETE firstname="Tiziana" nameprefix="" lastname="Papandrea" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:18:33.54">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Palermo" date="2023-05-21" nation="ITA" />
     <ATHLETE firstname="Tiziana" nameprefix="" lastname="Papandrea" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:31.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <ATHLETE firstname="Michelle" nameprefix="" lastname="Ware" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:07.87">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Crawley" date="2023-01-21" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:27.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Swansea" date="2020-02-29" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:34.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Riccione" date="2012-06-13" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:15.44">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2022-06-04" nation="GBR" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:44.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Aberdeen" date="2022-06-17" nation="GBR" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:29.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="2023-06-04" nation="GBR" />
     <ATHLETE firstname="Michelle" nameprefix="" lastname="Ware" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:07.55">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2022-09-04" nation="ITA" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:32.39">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Gwangju" date="2019-08-17" nation="KOR" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:33.61">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Aberdeen" date="2022-06-18" nation="GBR" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:05:32.44">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Riccione" date="2012-06-12" nation="ITA" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:27.09">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-06-28" nation="" />
     <ATHLETE firstname="Marie Therese" nameprefix="" lastname="Fuzzati" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:00.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-06" nation="" />
     <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:13.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-08-08" nation="" />
     <ATHLETE firstname="Jill" nameprefix="" lastname="Hernandez" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:40.66">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-08-11" nation="" />
     <ATHLETE firstname="Jill" nameprefix="" lastname="Hernandez" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:34.12">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-07-23" nation="" />
     <ATHLETE firstname="Susan" nameprefix="" lastname="Preston" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:18:15.80">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-07-29" nation="" />
     <ATHLETE firstname="Alison" nameprefix="" lastname="Zamanian" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:31.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-06-07" nation="" />
     <ATHLETE firstname="Cindy" nameprefix="" lastname="Mabee" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:07.87">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-01-21" nation="GBR" />
     <ATHLETE firstname="Joanna" nameprefix="" lastname="Corben" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:26.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2014-08-04" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:34.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Riccione" date="2012-06-13" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:15.44">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-06-04" nation="" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:44.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-06-17" nation="" />
     <ATHLETE firstname="Helen" nameprefix="" lastname="Gorman" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:29.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-07" nation="" />
     <ATHLETE firstname="Susan" nameprefix="" lastname="O'Neill" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:07.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2011-08-13" nation="" />
     <ATHLETE firstname="Jill" nameprefix="" lastname="Hernandez" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:31.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2001-08-18" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:31.02">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-08-07" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:20.68">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2014-08-05" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:29.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:01:05.73">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:02:28.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Cadiz" date="2009-09-16" nation="ESP" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:05:25.88">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Alkmaar" date="2018-04-08" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC Woerden" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:11:08.13">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Cadiz" date="2009-09-15" nation="ESP" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:21:31.80">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-04" nation="NED" />
     <ATHLETE firstname="Irene" nameprefix="van der" lastname="Laan" gender="F" nation="NED" CLUB="ZV De Bron" birthdate="1960-12-27" />
    </RECORD>
    <RECORD swimtime="00:00:35.46">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:01:17.35">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:02:46.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Cromjongh" gender="F" nation="NED" CLUB="De Zwoer" birthdate="1964-03-17" />
    </RECORD>
    <RECORD swimtime="00:00:38.31">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Ariene" nameprefix="" lastname="Knoester" gender="F" nation="NED" CLUB="Aqua-Novio&apos;94" birthdate="1967-09-28" />
    </RECORD>
    <RECORD swimtime="00:01:26.79">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Annette" nameprefix="" lastname="Wijnja-Visser" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1967-01-30" />
    </RECORD>
    <RECORD swimtime="00:03:06.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Annette" nameprefix="" lastname="Wijnja-Visser" gender="F" nation="NED" CLUB="De Biesboschzwemmers" birthdate="1967-01-30" />
    </RECORD>
    <RECORD swimtime="00:00:31.91">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1967-02-08" />
    </RECORD>
    <RECORD swimtime="00:01:16.54">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2013-09-03" nation="NED" />
     <ATHLETE firstname="Mathilde" nameprefix="" lastname="Vink" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1958-12-12" />
    </RECORD>
    <RECORD swimtime="00:03:00.68">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2013-09-04" nation="NED" />
     <ATHLETE firstname="Mathilde" nameprefix="" lastname="Vink" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1958-12-12" />
    </RECORD>
    <RECORD swimtime="00:02:48.67">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC Woerden" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:06:07.43">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Luxembourg" date="2018-10-13" nation="LUX" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC Woerden" birthdate="1963-05-15" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:28.84">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Fukuoka" date="2023-08-08" nation="JPN" />
     <ATHLETE firstname="Anette" nameprefix="" lastname="Philipsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:01:03.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gwangju" date="2019-08-13" nation="KOR" />
     <ATHLETE firstname="Susanne" nameprefix="" lastname="Reibel-Oberle" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:19.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Karlsruhe" date="2019-06-01" nation="GER" />
     <ATHLETE firstname="Susanne" nameprefix="" lastname="Reibel-Oberle" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:50.80">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gwangju" date="2019-08-18" nation="KOR" />
     <ATHLETE firstname="Susanne" nameprefix="" lastname="Reibel-Oberle" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:10:01.22">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Fukuoka" date="2023-08-05" nation="JPN" />
     <ATHLETE firstname="Claudia" nameprefix="" lastname="Thielemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:19:17.89">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Lodi" date="2022-06-11" nation="ITA" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Hoag" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:33.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Fukuoka" date="2023-08-11" nation="JPN" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:13.23">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Roma" date="2022-09-02" nation="ITA" />
     <ATHLETE firstname="Lise" nameprefix="" lastname="Lothe" gender="F" nation="NOR" />
    </RECORD>
    <RECORD swimtime="00:02:36.61">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Stratford" date="2019-03-24" nation="GBR" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Brown" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:35.94">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Treviso" date="2017-05-20" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:19.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Legnano" date="2017-01-29" nation="ITA" />
     <ATHLETE firstname="Pia" nameprefix="" lastname="Thulstrup" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:02:56.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Riccione" date="2019-12-08" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:30.65">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-07" nation="JPN" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:07.55">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-08" nation="JPN" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:36.33">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-10" nation="JPN" />
     <ATHLETE firstname="Claudia" nameprefix="" lastname="Thielemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:39.07">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gwangju" date="2019-08-15" nation="KOR" />
     <ATHLETE firstname="Susanne" nameprefix="" lastname="Reibel-Oberle" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:05:39.37">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gwangju" date="2019-08-14" nation="KOR" />
     <ATHLETE firstname="Susanne" nameprefix="" lastname="Reibel-Oberle" gender="F" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:27.94">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-04-21" nation="" />
     <ATHLETE firstname="Jennie" nameprefix="" lastname="Bucknell" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:01.87">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-04-20" nation="" />
     <ATHLETE firstname="Jennie" nameprefix="" lastname="Bucknell" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:02:16.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-08-06" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:43.41">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-07-10" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:09:44.76">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-02-25" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:18:36.30">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-07-08" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:31.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-08-02" nation="" />
     <ATHLETE firstname="Holly" nameprefix="" lastname="Geen Blair" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:09.69">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-11-08" nation="" />
     <ATHLETE firstname="Holly" nameprefix="" lastname="Geen Blair" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:31.79">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-05-19" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:35.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-08-11" nation="" />
     <ATHLETE firstname="Andrea" nameprefix="" lastname="Muller" gender="F" nation="CHI" />
    </RECORD>
    <RECORD swimtime="00:01:19.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-01-29" nation="" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:57.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-08-10" nation="" />
     <ATHLETE firstname="Andrea" nameprefix="" lastname="Muller" gender="F" nation="CHI" />
    </RECORD>
    <RECORD swimtime="00:00:30.43">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-07" nation="" />
     <ATHLETE firstname="Andrea" nameprefix="" lastname="Muller" gender="F" nation="CHI" />
    </RECORD>
    <RECORD swimtime="00:01:07.55">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-08" nation="" />
     <ATHLETE firstname="Franca" nameprefix="" lastname="Bosisio" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:36.33">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-10" nation="" />
     <ATHLETE firstname="Claudia" nameprefix="" lastname="Thielemann" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:31.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-06-07" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:22.41">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-06-07" nation="" />
     <ATHLETE firstname="Ellen" nameprefix="" lastname="Reynolds" gender="F" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:30.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:01:08.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-15" nation="HUN" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:02:33.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Londen" date="2016-05-26" nation="GBR" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:05:26.24">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg" date="2017-10-14" nation="LUX" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:11:26.49">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2012-06-10" nation="ITA" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:22:17.27">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-02" nation="NED" />
     <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" CLUB="PSV" birthdate="1959-04-01" />
    </RECORD>
    <RECORD swimtime="00:00:37.72">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Londen" date="2016-05-27" nation="GBR" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:01:24.02">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:03:00.41">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Luxembourg" date="2016-10-15" nation="LUX" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:00:43.06">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Linda" nameprefix="van de" lastname="Ree" gender="F" nation="NED" CLUB="De Ganze" birthdate="1963-10-26" />
    </RECORD>
    <RECORD swimtime="00:01:32.45">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-09-04" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:03:28.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Montreal" date="2014-08-08" nation="CAN" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:00:34.14">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:01:21.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:03:18.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Margriet" nameprefix="" lastname="Grove-Lingeman" gender="F" nation="NED" CLUB="Triton" birthdate="1962-02-05" />
    </RECORD>
    <RECORD swimtime="00:02:52.46">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-05-15" />
    </RECORD>
    <RECORD swimtime="00:06:40.81">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" CLUB="PSV" birthdate="1959-04-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:29.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <ATHLETE firstname="Dawn" nameprefix="" lastname="Kissack" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:06.02">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Madrid" date="2021-06-13" nation="ESP" />
     <ATHLETE firstname="Carmen" nameprefix="" lastname="Navarro" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:27.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="Carmen" nameprefix="" lastname="Navarro" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:05:15.75">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2022-08-29" nation="ITA" />
     <ATHLETE firstname="Barbara" nameprefix="" lastname="Gellrich" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:10:58.35">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2016-06-21" nation="ITA" />
     <ATHLETE firstname="Cristina" nameprefix="" lastname="Tarantino" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:21:12.79">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-04" nation="GBR" />
     <ATHLETE firstname="Suzanne" nameprefix="" lastname="Noble" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:35.09">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <ATHLETE firstname="Julie" nameprefix="" lastname="Hoyle" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:16.63">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Aberdeen" date="2022-06-19" nation="GBR" />
     <ATHLETE firstname="Julie" nameprefix="" lastname="Hoyle" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:46.79">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Aberdeen" date="2022-06-18" nation="GBR" />
     <ATHLETE firstname="Julie" nameprefix="" lastname="Hoyle" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:37.43">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Lignano" date="2022-02-06" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:23.04">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Trevisio" date="2022-05-20" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:03:06.40">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2022-09-01" nation="ITA" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:32.36">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Madrid" date="2022-06-19" nation="ESP" />
     <ATHLETE firstname="Carmen" nameprefix="" lastname="Navarro" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:14.21">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Las Palmas" date="2022-07-11" nation="ESP" />
     <ATHLETE firstname="Carmen" nameprefix="" lastname="Navarro" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:49.71">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Lodi" date="2023-06-11" nation="ITA" />
     <ATHLETE firstname="Daniela" nameprefix="" lastname="Pedacchiola" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:48.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="London" date="2016-05-25" nation="GBR" />
     <ATHLETE firstname="Colette" nameprefix="" lastname="Crabbe" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:01.90">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <ATHLETE firstname="Colette" nameprefix="" lastname="Crabbe" gender="F" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:28.84">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-05" nation="" />
     <ATHLETE firstname="Holly" nameprefix="" lastname="Green" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:03.83">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2011-08-05" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:21.03">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-03-20" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:04:53.58">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-06-11" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:10:06.23">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-02-11" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:19:23.70">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-06-18" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:00:33.38">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-08-05" nation="" />
     <ATHLETE firstname="Holly" nameprefix="" lastname="Green" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:14.28">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-08-13" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:41.38">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-05-13" nation="" />
     <ATHLETE firstname="Karlyn" nameprefix="" lastname="Pipes-Neilsen" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:37.43">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-02-06" nation="" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:23.07">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-02-06" nation="" />
     <ATHLETE firstname="Monica" nameprefix="" lastname="Coro" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:03:04.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-03-18" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:00:29.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-04" nation="" />
     <ATHLETE firstname="Holly" nameprefix="" lastname="Green" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:12.06">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2011-08-04" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:41.03">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2011-08-06" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:44.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-03-20" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:05:48.88">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-06-11" nation="" />
     <ATHLETE firstname="Lynn" nameprefix="" lastname="Marshall" gender="F" nation="CAN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:31.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:01:09.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:02:37.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rome" date="2022-08-31" nation="ITA" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:05:39.78">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Alkmaar" date="2022-04-10" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:11:47.84">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:22:41.46">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg" date="2019-10-12" nation="LUX" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:00:38.83">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:01:22.93">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:02:59.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rome" date="2022-09-01" nation="ITA" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:00:44.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:01:35.58">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kranj" date="2018-09-07" nation="SLO" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:03:27.58">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kranj" date="2018-09-04" nation="SLO" />
     <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" CLUB="PSV" birthdate="1953-04-03" />
    </RECORD>
    <RECORD swimtime="00:00:36.68">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2017-05-06" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:01:34.35">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Luxembourg/Hollerich" date="2022-10-08" nation="LUX" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:04:23.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Nijmegen" date="2000-06-10" nation="NED" />
     <ATHLETE firstname="Annie" nameprefix="de" lastname="Vos" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1934-01-10" />
    </RECORD>
    <RECORD swimtime="00:03:09.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Luxembourg/Hollerich" date="2021-10-10" nation="LUX" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
    <RECORD swimtime="00:07:05.68">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Luxembourg/Hollerich" date="2022-10-08" nation="LUX" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1956-12-31" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:30.56">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <ATHLETE firstname="Alyson" nameprefix="" lastname="Fordham" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:09.16">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-04" nation="GBR" />
     <ATHLETE firstname="Alyson" nameprefix="" lastname="Fordham" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:37.34">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rome" date="2022-08-31" nation="ITA" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:05:33.65">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Citavecchia" date="2021-06-29" nation="ITA" />
     <ATHLETE firstname="Cristina" nameprefix="" lastname="Tarantino" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:11:32.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Civitavecchia" date="2021-06-29" nation="ITA" />
     <ATHLETE firstname="Cristina" nameprefix="" lastname="Tarantino" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:21:56.07">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Glasgow" date="2019-11-09" nation="GBR" />
     <ATHLETE firstname="Audrey" nameprefix="" lastname="Cooper" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:37.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Yalta" date="2011-09-07" nation="UKR" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:01:21.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="G�teborg" date="2010-08-05" nation="SWE" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:02:59.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rome" date="2022-09-01" nation="ITA" />
     <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:40.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Braunschweig" date="2021-09-11" nation="GER" />
     <ATHLETE firstname="Dagmar" nameprefix="" lastname="Frese" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:29.97">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <ATHLETE firstname="Esther" nameprefix="" lastname="Iseppi" gender="F" nation="SUI" />
    </RECORD>
    <RECORD swimtime="00:03:12.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Aberdeen" date="2022-06-17" nation="GBR" />
     <ATHLETE firstname="Amanda" nameprefix="" lastname="Heath" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:35.27">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Aberdeen" date="2022-06-18" nation="GBR" />
     <ATHLETE firstname="Lindsey" nameprefix="" lastname="Gowland" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:20.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Colette" nameprefix="" lastname="Crabbe" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:03:16.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <ATHLETE firstname="Amanda" nameprefix="" lastname="Heath" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:55.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Colette" nameprefix="" lastname="Crabb�" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:06:21.10">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Colette" nameprefix="" lastname="Crabb�" gender="F" nation="BEL" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:29.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-03-08" nation="" />
     <ATHLETE firstname="Penny" nameprefix="" lastname="Noyes" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:04.89">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-07-30" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:25.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-08-18" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:12.80">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-10-08" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:10:49.60">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-07-15" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:20:41.53">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-07-21" nation="" />
     <ATHLETE firstname="S." nameprefix="" lastname="Heim-Bowen" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:33.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-08-02" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:14.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-07-31" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:47.70">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-08-08" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:39.91">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-04-02" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:28.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-05-25" nation="" />
     <ATHLETE firstname="Jenny" nameprefix="" lastname="Whiteley" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:03:12.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-06-17" nation="" />
     <ATHLETE firstname="Amanda" nameprefix="" lastname="Heath" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:32.36">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-07" nation="" />
     <ATHLETE firstname="Traci" nameprefix="" lastname="Granger" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:13.70">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2016-08-18" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:57.26">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-07-20" nation="" />
     <ATHLETE firstname="Penny" nameprefix="" lastname="Noyes" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:51.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-04-08" nation="" />
     <ATHLETE firstname="Penny" nameprefix="" lastname="Noyes" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:14.58">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-07-19" nation="" />
     <ATHLETE firstname="Penny" nameprefix="" lastname="Noyes" gender="F" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:33.80">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:01:16.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:01:16.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Rome" date="2022-09-04" nation="ITA" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="SWOL1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:02:56.90">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:06:38.57">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg/Hollerich" date="2021-10-09" nation="LUX" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:13:29.34">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg/Hollerich" date="2021-10-09" nation="LUX" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:25:25.33">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg/Hollerich" date="2021-10-09" nation="LUX" />
     <ATHLETE firstname="Conny" nameprefix="" lastname="Boer-Buijs" gender="F" nation="NED" CLUB="ZVVS" birthdate="1950-11-30" />
    </RECORD>
    <RECORD swimtime="00:00:44.81">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Oosterhout" date="2017-04-09" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:01:41.30">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Luxembourg" date="2016-10-16" nation="LUX" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:03:45.13">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:00:46.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:01:48.98">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Oosterhout" date="2016-04-10" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:03:58.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Luxembourg" date="2017-10-14" nation="LUX" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:00:40.27">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:01:44.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:04:50.47">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Halle" date="2004-08-16" nation="GER" />
     <ATHLETE firstname="Annie" nameprefix="de" lastname="Vos" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1934-01-10" />
    </RECORD>
    <RECORD swimtime="00:03:27.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" CLUB="Swol 1894" birthdate="1951-05-17" />
    </RECORD>
    <RECORD swimtime="00:08:51.69">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Halle" date="2004-08-16" nation="GER" />
     <ATHLETE firstname="Annie" nameprefix="de" lastname="Vos" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1934-01-10" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:32.63">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2023-05-14" nation="ITA" />
     <ATHLETE firstname="Carole Wendy" nameprefix="" lastname="Smith" gender="F" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:15.01">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gera" date="2010-03-13" nation="GER" />
     <ATHLETE firstname="Christel" nameprefix="" lastname="Schulz" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:48.03">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="G�teborg" date="2010-08-02" nation="SWE" />
     <ATHLETE firstname="Christel" nameprefix="" lastname="Schulz" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:06:04.56">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Mulhouse" date="2022-06-25" nation="FRA" />
     <ATHLETE firstname="Martine" nameprefix="" lastname="Reynaud" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:12:32.21">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Christchurch" date="2002-03-24" nation="NZL" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:24:06.48">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Glasgow" date="2001-06-01" nation="SCO" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:38.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Turku" date="2015-10-24" nation="FIN" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:01:25.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:03:06.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Turku" date="2015-10-24" nation="FIN" />
     <ATHLETE firstname="Margit" nameprefix="" lastname="Ohlsson" gender="F" nation="SWE" />
    </RECORD>
    <RECORD swimtime="00:00:41.67">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Hannover" date="2014-06-22" nation="GER" />
     <ATHLETE firstname="Monika" nameprefix="" lastname="Senftleben" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:37.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Swansea" date="2013-03-09" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:30.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Plymouth" date="2013-06-14" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:36.36">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Montreal" date="2014-08-05" nation="CAN" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:24.55">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Montreal" date="2014-08-06" nation="CAN" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:40.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Montreal" date="2014-08-08" nation="CAN" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:10.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="London" date="2016-05-25" nation="GBR" />
     <ATHLETE firstname="Brigitte" nameprefix="" lastname="Merten" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:06:54.30">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Berlin" date="2016-01-23" nation="GER" />
     <ATHLETE firstname="Brigitte" nameprefix="" lastname="Merten" gender="F" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:30.73">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-09" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:06.68">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-06" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:29.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-14" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:21.19">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-13" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:11:04.90">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-06-03" nation="" />
     <ATHLETE firstname="Christie" nameprefix="" lastname="Ciraulo" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:21:02.79">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-02" nation="" />
     <ATHLETE firstname="Christie" nameprefix="" lastname="Ciraulo" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:34.65">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-10" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:16.27">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-08-04" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:49.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-08" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:41.67">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Hannover" date="2014-06-22" nation="GER" />
     <ATHLETE firstname="Monika" nameprefix="" lastname="Senftleben" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:35.93">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-10-02" nation="" />
     <ATHLETE firstname="Nobuko" nameprefix="" lastname="Yasuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:29.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-07-15" nation="" />
     <ATHLETE firstname="Nobuko" nameprefix="" lastname="Yasuda" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:34.68">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-07-23" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:16.07">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-10-08" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:21.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-05-27" nation="" />
     <ATHLETE firstname="Andra" nameprefix="" lastname="Jaunzeme" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:00.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-08-01" nation="USA" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:45.75">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-05-28" nation="" />
     <ATHLETE firstname="Laura" nameprefix="" lastname="Vaca" gender="F" nation="MEX" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:37.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:01:28.01">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2021-09-12" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:03:15.74">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="G�teborg" date="2010-08-02" nation="SWE" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:07:04.33">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="G�teborg" date="2010-08-06" nation="SWE" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:14:59.75">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="G�teborg" date="2010-07-31" nation="SWE" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:28:55.03">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-05" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:00:51.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2012-05-06" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:55.72">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2011-05-06" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:04:12.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2010-05-07" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:00:48.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Rome" date="2022-09-02" nation="ITA" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:01:52.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="00:04:26.89">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kampen" date="2004-04-24" nation="NED" />
     <ATHLETE firstname="Ati" nameprefix="" lastname="Derkse-den Boer" gender="F" nation="NED" CLUB="Aquapoldro" birthdate="1929-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:55.26">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Luxembourg/Hollerich" date="2021-10-10" nation="LUX" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:03:49.47">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Luxembourg/Hollerich" date="2021-10-10" nation="LUX" />
     <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" CLUB="PSV" birthdate="1946-12-26" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:34.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2006-03-03" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:20.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kazan" date="2015-08-11" nation="RUS" />
     <ATHLETE firstname="Christel" nameprefix="" lastname="Schulz" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:56.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Perth" date="2008-04-20" nation="AUS" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:06:13.20">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="San Francisco" date="2006-08-10" nation="USA" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:12:58.94">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg" date="2006-10-22" nation="LUX" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:24:41.76">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2006-03-03" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:42.72">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Hillerod" date="2018-06-16" nation="DEN" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:01:33.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Hillerod" date="2018-06-16" nation="DEN" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:03:23.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Hillerod" date="2018-06-17" nation="DEN" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:00:46.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Cadiz" date="2009-09-16" nation="ESP" />
     <ATHLETE firstname="Eliane" nameprefix="" lastname="Pellis" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:01:42.27">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Swansea" date="2019-06-15" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:43.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Gera" date="2014-04-04" nation="GER" />
     <ATHLETE firstname="Luise" nameprefix="" lastname="Kn�pfle" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:38.93">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Vichy" date="2019-05-25" nation="FRA" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:34.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Chalon" date="2019-06-23" nation="FRA" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:04:03.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Riccione" date="2004-06-09" nation="ITA" />
     <ATHLETE firstname="Sylvia" nameprefix="" lastname="Neuhauser" gender="F" nation="AUT" />
    </RECORD>
    <RECORD swimtime="00:03:21.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Braunschweig" date="2022-04-22" nation="GER" />
     <ATHLETE firstname="Kira" nameprefix="" lastname="Makarova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:07:29.06">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Roma" date="2022-08-30" nation="ITA" />
     <ATHLETE firstname="Brigitte" nameprefix="" lastname="Merten" gender="F" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:34.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-08" nation="" />
     <ATHLETE firstname="Diann" nameprefix="" lastname="Uustal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:17.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-09" nation="" />
     <ATHLETE firstname="Diann" nameprefix="" lastname="Uustal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:54.26">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-09-27" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:06:12.25">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-07-12" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:12:58.94">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg" date="2006-10-22" nation="LUX" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:24:41.76">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2006-03-03" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:40.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-09" nation="" />
     <ATHLETE firstname="Diann" nameprefix="" lastname="Uustal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:28.67">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-10-10" nation="" />
     <ATHLETE firstname="Diann" nameprefix="" lastname="Uustal" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:16.80">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-04-28" nation="" />
     <ATHLETE firstname="Clary" nameprefix="" lastname="Munns" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:00:43.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-03-06" nation="" />
     <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:38.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-03-06" nation="" />
     <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:40.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2014-07-19" nation="" />
     <ATHLETE firstname="Joann" nameprefix="" lastname="Leilich" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:38.93">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-05-25" nation="" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:34.88">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-06-23" nation="" />
     <ATHLETE firstname="Judith" nameprefix="" lastname="Wilson" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:44.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-04-28" nation="" />
     <ATHLETE firstname="Clary" nameprefix="" lastname="Munns" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:03:21.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-04-22" nation="" />
     <ATHLETE firstname="Kira" nameprefix="" lastname="Makarova" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:07:39.96">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Swansea" date="2006-03-03" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:40.60">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-07" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:34.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-15" nation="HUN" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:03:40.81">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-16" nation="HUN" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:07:56.27">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:16:15.33">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2015-05-08" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:31:22.53">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg" date="2017-10-14" nation="LUX" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:00:54.51">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" CLUB="PSV" birthdate="1935-10-12" />
    </RECORD>
    <RECORD swimtime="00:02:02.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2015-05-10" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:04:28.02">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2015-05-10" nation="NED" />
     <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" CLUB="PSV" birthdate="1935-10-12" />
    </RECORD>
    <RECORD swimtime="00:01:06.15">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sydney" date="2009-10-15" nation="AUS" />
     <ATHLETE firstname="Anneke" nameprefix="" lastname="Logtenberg" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1929-10-31" />
    </RECORD>
    <RECORD swimtime="00:02:25.55">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Luxembourg" date="2017-10-15" nation="LUX" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:05:28.40">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sydney" date="2009-10-16" nation="AUS" />
     <ATHLETE firstname="Anneke" nameprefix="" lastname="Logtenberg" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1929-10-31" />
    </RECORD>
    <RECORD swimtime="00:01:07.79">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:02:29.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:37.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Leeds" date="2011-06-18" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:24.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Leeds" date="2011-06-19" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:07.40">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2011-03-06" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:06:39.90">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2012-05-05" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:13:51.21">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Crawley" date="2011-01-29" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:26:29.87">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2011-03-04" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:46.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Fukuoka" date="2023-08-11" nation="JPN" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:01:39.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Gentofte" date="2023-05-29" nation="DEN" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:03:41.85">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Solingen" date="2022-03-19" nation="GER" />
     <ATHLETE firstname="Christel" nameprefix="" lastname="Schulz" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:46.94">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2023-06-02" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:43.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:51.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Sheffield" date="2023-06-04" nation="GBR" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:46.21">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Leeds" date="2011-06-17" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:01.54">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Cadiz" date="2009-09-16" nation="ESP" />
     <ATHLETE firstname="Sylvia" nameprefix="" lastname="Neuhauser" gender="F" nation="AUT" />
    </RECORD>
    <RECORD swimtime="00:04:22.67">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Cadiz" date="2009-09-17" nation="ESP" />
     <ATHLETE firstname="Sylvia" nameprefix="" lastname="Neuhauser" gender="F" nation="AUT" />
    </RECORD>
    <RECORD swimtime="00:03:54.07">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Cardiff" date="2011-05-06" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:21.88">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Crawley" date="2011-01-30" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:36.61">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-07-15" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:23.16">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-07-14" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:05.95">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-09-20" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:06:39.90">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2012-05-05" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:13:51.21">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Crawley" date="2011-01-29" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:28:35.98">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-03-11" nation="" />
     <ATHLETE firstname="Denise" nameprefix="" lastname="Robertson" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:00:43.04">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-03-11" nation="" />
     <ATHLETE firstname="Satoko" nameprefix="" lastname="Takeuji" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:39.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-05-29" nation="" />
     <ATHLETE firstname="Elisabeth" nameprefix="" lastname="Ketelsen" gender="F" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:03:32.61">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-06-04" nation="" />
     <ATHLETE firstname="Noriko" nameprefix="" lastname="Yoshida" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:46.94">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-06-02" nation="" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:43.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-06-03" nation="" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:51.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-06-04" nation="" />
     <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:46.21">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Leeds" date="2011-06-17" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:54.93">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2012-04-21" nation="" />
     <ATHLETE firstname="Judie" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:04:15.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2012-07-14" nation="" />
     <ATHLETE firstname="Judie" nameprefix="" lastname="Oliver" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:03:53.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-08-17" nation="" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:08:21.88">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Crawley" date="2011-01-30" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:48.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:55.92">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg/Hollerich" date="2022-10-08" nation="LUX" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:04:14.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg/Hollerich" date="2021-10-10" nation="LUX" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:08:56.64">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2021-09-12" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:18:55.00">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-05" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:35:55.82">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-05" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:01.74">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:02:19.73">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rome" date="2022-09-02" nation="ITA" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:05:02.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Luxembourg/Hollerich" date="2022-10-08" nation="LUX" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:29.00">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2012-05-05" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:02:58.82">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Luxembourg/Hollerich" date="2021-10-10" nation="LUX" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:06:45.88">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2021-09-12" nation="NED" />
     <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" CLUB="PSV" birthdate="1935-09-21" />
    </RECORD>
    <RECORD swimtime="00:01:11.26">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="00:02:29.94">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Marie" nameprefix="" lastname="Smits" gender="F" nation="NED" CLUB="Old Dutch" birthdate="1938-12-30" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:38.98">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2016-05-27" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:29.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Norwich" date="2016-05-07" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:31.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2016-05-26" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:07:03.60">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg" date="2016-10-15" nation="LUX" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:14:27.71">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2016-04-01" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:28:11.18">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2016-03-05" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:48.85">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Gyula" date="2019-06-29" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:01:45.27">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Gyula" date="2019-06-30" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:03:43.27">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Gyula" date="2019-06-28" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:00:51.83">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:01:54.96">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:04:18.23">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:00:48.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Gwangju" date="2019-08-14" nation="KOR" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:04.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Gyula" date="2019-06-29" nation="HUN" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:06:18.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Schiltighem" date="2016-05-08" nation="FRA" />
     <ATHLETE firstname="Yvette" nameprefix="" lastname="Kaplan Bader" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:03:54.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gwangju" date="2019-08-15" nation="KOR" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:11:16.32">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Millau" date="2014-07-05" nation="FRA" />
     <ATHLETE firstname="Yvette" nameprefix="" lastname="Kaplan Bader" gender="F" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:38.89">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-08" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:27.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-06" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:14.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-07" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:07:03.60">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-10-15" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:14:27.71">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-04-01" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:28:11.18">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-03-05" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:47.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-09-18" nation="" />
     <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:45.27">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-06-30" nation="" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:03:43.27">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-08-13" nation="" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:00:51.83">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:01:54.96">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:04:18.23">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:00:48.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-08-14" nation="" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:01.26">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-09-11" nation="" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:05:07.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2009-07-25" nation="" />
     <ATHLETE firstname="Lois Kivi" nameprefix="" lastname="Nochman" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:54.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-08-15" nation="" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:08:26.93">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-09-11" nation="" />
     <ATHLETE firstname="Katharina" nameprefix="" lastname="Flora" gender="F" nation="HUN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:01:16.67">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:14.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-07" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:07:15.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:31.61">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2017-05-05" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:19.12">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2016-05-07" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:06:55.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2016-05-07" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:01:43.32">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Oosterhout" date="2017-04-09" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:46.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:08:13.89">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:00:45.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Crawley" date="2022-01-23" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:46.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Aberdeen" date="2022-06-18" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:52.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Aberdeen" date="2022-06-19" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:25.92">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2022-03-05" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:18:18.20">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:34:29.59">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:54.49">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Crawley" date="2022-01-23" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:59.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Crawley" date="2022-01-23" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:04:32.59">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Crawley" date="2022-01-23" nation="GBR" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:59.40">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kortrijk" date="2023-11-05" nation="BEL" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:02:14.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kortrijk" date="2023-11-04" nation="BEL" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:04:53.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Charleroi" date="2022-11-02" nation="BEL" />
     <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:00:45.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-01-23" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:46.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-06-18" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:52.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-06-19" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:08:25.92">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-03-05" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:18:18.20">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-09-11" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:33:36.10">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2020-02-21" nation="" />
     <ATHLETE firstname="Dorothy" nameprefix="" lastname="Dickey" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:00:54.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-01-23" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:59.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-01-23" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:04:32.89">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-01-23" nation="" />
     <ATHLETE firstname="Jane" nameprefix="" lastname="Asher" gender="F" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:03.72">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-09-03" nation="NED" />
     <ATHLETE firstname="Olga" nameprefix="" lastname="Kokorina" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:27.19">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2013-06-02" nation="" />
     <ATHLETE firstname="Olga" nameprefix="" lastname="Kokorina" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:05:21.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2013-06-01" nation="RUS" />
     <ATHLETE firstname="Olga" nameprefix="" lastname="Kokorina" gender="F" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:22.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2012-07-16" nation="" />
     <ATHLETE firstname="Yone" nameprefix="" lastname="Murata" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:39.01">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2014-08-06" nation="" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Ronai" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:08:52.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2014-08-08" nation="" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Ronai" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:06:30.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2008-08-16" nation="" />
     <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:14:12.52">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2014-08-05" nation="" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Ronai" gender="F" nation="BRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:01:21.48">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2021-09-12" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:56.62">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:43.62">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:03:43.56">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:07.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:04:35.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="00:09:51.05">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2021-09-12" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" CLUB="PSV" birthdate="1926-10-08" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:01:07.27">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kaerepere" date="2017-02-04" nation="EST" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Kutti" gender="F" nation="EST" />
    </RECORD>
    <RECORD swimtime="00:03:56.62">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:08:57.23">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="St. Germain" date="2006-03-25" nation="FRA" />
     <ATHLETE firstname="Marie" nameprefix="de" lastname="Fromont" gender="F" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:18:16.28">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Barcelona" date="2007-05-26" nation="ESP" />
     <ATHLETE firstname="Bernarda" nameprefix="" lastname="Angulo" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="00:01:30.96">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Gera" date="2016-04-17" nation="GER" />
     <ATHLETE firstname="Ingeborg" nameprefix="" lastname="Fritze" gender="F" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:43.56">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:08:49.98">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Madrid" date="2009-07-31" nation="ESP" />
     <ATHLETE firstname="Bernarda" nameprefix="" lastname="Angulo" gender="F" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:07.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:04:35.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:09:51.05">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2021-09-12" nation="NED" />
     <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:01:03.25">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-04-02" nation="" />
     <ATHLETE firstname="Liz" nameprefix="" lastname="Wallis" gender="F" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:02:22.74">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-08-07" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:03.47">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-08-18" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:10:12.49">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-08-06" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:21:39.10">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-14" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:41:39.68">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-06-02" nation="" />
     <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:14.31">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2013-08-10" nation="" />
     <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:42.67">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2013-08-08" nation="" />
     <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:42.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2016-05-29" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:38.21">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-06-23" nation="" />
     <ATHLETE firstname="Kalis" nameprefix="" lastname="Rasmussen" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:03:23.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-09-17" nation="" />
     <ATHLETE firstname="Teruko" nameprefix="" lastname="Ono" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:07:42.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-06-23" nation="" />
     <ATHLETE firstname="Kalis" nameprefix="" lastname="Rasmussen" gender="F" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:56.76">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-04-14" nation="" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Ronai" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:05:12.53">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-12-04" nation="" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Ronai" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:12:05.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-11-16" nation="" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Ronai" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:08:51.10">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-11-15" nation="" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Ronai" gender="F" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:18:50.06">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-11-04" nation="" />
     <ATHLETE firstname="Nora" nameprefix="" lastname="Ronai" gender="F" nation="BRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="00:01:12.84">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-07-31" nation="USA" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:52.45">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-07-11" nation="" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:33.32">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-07-31" nation="USA" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:16:36.80">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-01-19" nation="" />
     <ATHLETE firstname="Mieko" nameprefix="" lastname="Nagaoka" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:38:04.30">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-06-15" nation="" />
     <ATHLETE firstname="Mieko" nameprefix="" lastname="Nagaoka" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="01:14:08.73">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-06-14" nation="" />
     <ATHLETE firstname="Mieko" nameprefix="" lastname="Nagaoka" gender="F" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:29.84">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-08-01" nation="USA" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:04.26">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-07-31" nation="USA" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:40.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-07-11" nation="USA" />
     <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="20" agemax="24" />
   <RECORDS>
    <RECORD swimtime="00:00:23.24">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Brandon" nameprefix="van den" lastname="Berg" gender="M" nation="NED" CLUB="Blue Marlins (SG)" birthdate="2002-05-23" />
    </RECORD>
    <RECORD swimtime="00:00:51.62">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Brandon" nameprefix="van den" lastname="Berg" gender="M" nation="NED" CLUB="Blue Marlins (SG)" birthdate="2002-05-23" />
    </RECORD>
    <RECORD swimtime="00:01:54.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Maquinho" nameprefix="" lastname="Vorst" gender="M" nation="NED" CLUB="De Dinkel" birthdate="2002-03-04" />
    </RECORD>
    <RECORD swimtime="00:04:17.05">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="startlimiet" nameprefix="" lastname="" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:08:59.66">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="startlimiet" nameprefix="" lastname="" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:17:10.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-04" nation="NED" />
     <ATHLETE firstname="Janne" nameprefix="" lastname="Englebert" gender="M" nation="NED" CLUB="Hieronymus" birthdate="2001-03-04" />
    </RECORD>
    <RECORD swimtime="00:00:26.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:00:57.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:02:10.58">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2014-05-04" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Albion" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:00:29.53">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <ATHLETE firstname="Coen" nameprefix="de" lastname="Bruijn" gender="M" nation="NED" CLUB="Hieronymus" birthdate="1992-07-06" />
    </RECORD>
    <RECORD swimtime="00:01:05.14">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2015-05-08" nation="NED" />
     <ATHLETE firstname="Coen" nameprefix="de" lastname="Bruijn" gender="M" nation="NED" CLUB="Hieronymus" birthdate="1992-07-06" />
    </RECORD>
    <RECORD swimtime="00:02:25.31">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Den Haag" date="2014-05-03" nation="NED" />
     <ATHLETE firstname="Roald" nameprefix="" lastname="Blok" gender="M" nation="NED" CLUB="Octopus" birthdate="1993-01-06" />
    </RECORD>
    <RECORD swimtime="00:00:25.06">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2015-05-08" nation="NED" />
     <ATHLETE firstname="Sverre" nameprefix="" lastname="Eschweiler" gender="M" nation="NED" CLUB="De Golfbreker" birthdate="1992-11-17" />
    </RECORD>
    <RECORD swimtime="00:00:56.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:02:05.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Albion" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:02:10.80">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2014-05-02" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Albion" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:04:51.88">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Nicko" nameprefix="" lastname="Kamphuis" gender="M" nation="NED" CLUB="De Warande" birthdate="1999-07-08" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:23.38">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Feijenoord Zwemmen (SG)" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:00:51.37">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-05-10" nation="NED" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Oosting" gender="M" nation="NED" CLUB="PSV" birthdate="1981-04-01" />
    </RECORD>
    <RECORD swimtime="00:01:54.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-05-10" nation="NED" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Oosting" gender="M" nation="NED" CLUB="PSV" birthdate="1981-04-01" />
    </RECORD>
    <RECORD swimtime="00:04:12.70">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-05-09" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:08:41.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-05-09" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:16:44.41">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-05-08" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:00:26.75">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Feijenoord Albion zwemclub" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:00:57.51">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" CLUB="Feijenoord Albion zwemclub" birthdate="1994-02-18" />
    </RECORD>
    <RECORD swimtime="00:02:13.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Riccione" date="2004-06-06" nation="ITA" />
     <ATHLETE firstname="Dennis" nameprefix="" lastname="Brouwers" gender="M" nation="NED" CLUB="Njord" birthdate="1978-07-14" />
    </RECORD>
    <RECORD swimtime="00:00:29.16">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2011-05-07" nation="NED" />
     <ATHLETE firstname="Rudy Ted" nameprefix="de" lastname="Haan" gender="M" nation="NED" CLUB="Anker Team Groningen" birthdate="1984-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:04.61">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2009-05-10" nation="NED" />
     <ATHLETE firstname="Rudy Ted" nameprefix="de" lastname="Haan" gender="M" nation="NED" CLUB="Anker Team Groningen" birthdate="1984-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:25.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Den Haag" date="2014-05-03" nation="NED" />
     <ATHLETE firstname="Tim" nameprefix="van den" lastname="Berg" gender="M" nation="NED" CLUB="MNC Dordrecht" birthdate="1985-04-13" />
    </RECORD>
    <RECORD swimtime="00:00:23.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Verhoeven" gender="M" nation="NED" CLUB="Feijenoord Albion zwemclub" birthdate="1997-04-18" />
    </RECORD>
    <RECORD swimtime="00:00:57.06">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2014-05-02" nation="NED" />
     <ATHLETE firstname="Filipp" nameprefix="" lastname="M�ller" gender="M" nation="NED" CLUB="Piranha" birthdate="1986-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:12.82">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2008-01-19" nation="NED" />
     <ATHLETE firstname="Rory Bob" nameprefix="de" lastname="Haan" gender="M" nation="NED" CLUB="Anker Team Groningen" birthdate="1981-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:12.58">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2011-05-07" nation="NED" />
     <ATHLETE firstname="Raymond" nameprefix="van der" lastname="Merwe" gender="M" nation="NED" CLUB="WVZ" birthdate="1986-11-19" />
    </RECORD>
    <RECORD swimtime="00:04:42.78">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2011-05-08" nation="NED" />
     <ATHLETE firstname="Raymond" nameprefix="van der" lastname="Merwe" gender="M" nation="NED" CLUB="WVZ" birthdate="1986-11-19" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:22.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Jyv�skyl�" date="2017-02-18" nation="FIN" />
     <ATHLETE firstname="Ari-Pekka" nameprefix="" lastname="Liukkonen" gender="M" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:00:50.81">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Aalto Alvari" date="2014-10-26" nation="FIN" />
     <ATHLETE firstname="Ari-Pekka" nameprefix="" lastname="Liukkonen" gender="M" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:01:50.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-16" nation="HUN" />
     <ATHLETE firstname="David" nameprefix="" lastname="Alcolado" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:04:00.96">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Palma de Mallorca" date="2022-06-05" nation="ESP" />
     <ATHLETE firstname="Alexander" nameprefix="" lastname="Fedorov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:08:27.48">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-12" nation="GER" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Dmitriev" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:16:13.78">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Barcelona" date="2015-04-12" nation="ESP" />
     <ATHLETE firstname="Rafael" nameprefix="" lastname="Cabanillas" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:25.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Penza" date="2016-04-03" nation="RUS" />
     <ATHLETE firstname="Anton" nameprefix="" lastname="Butymov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:56.20">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kazan" date="2015-08-15" nation="RUS" />
     <ATHLETE firstname="Vitalij" nameprefix="" lastname="Borisov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:02.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Obninsk" date="2019-04-26" nation="RUS" />
     <ATHLETE firstname="Dmitri" nameprefix="" lastname="Gorbunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:27.21">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Saransk" date="2021-04-18" nation="RUS" />
     <ATHLETE firstname="Kirill" nameprefix="" lastname="Strelnikov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:00.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Saransk" date="2021-04-16" nation="RUS" />
     <ATHLETE firstname="Kirill" nameprefix="" lastname="Strelnikov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:17.51">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Linz" date="2018-10-26" nation="AUT" />
     <ATHLETE firstname="Johannes" nameprefix="" lastname="Dietrich" gender="M" nation="AUT" />
    </RECORD>
    <RECORD swimtime="00:00:23.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Verhoeven" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:00:54.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Swansea" date="2008-03-02" nation="GBR" />
     <ATHLETE firstname="Matthew" nameprefix="" lastname="Bowe" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:00.74">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="St. Petersburg" date="2022-06-05" nation="RUS" />
     <ATHLETE firstname="Aleksandr" nameprefix="" lastname="Pribytok" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:03.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Obninsk" date="2019-04-28" nation="RUS" />
     <ATHLETE firstname="Dmitri" nameprefix="" lastname="Gorbunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:04:31.47">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Montreal" date="1994-07-06" nation="CAN" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="25" agemax="29" />
   <RECORDS>
    <RECORD swimtime="00:00:22.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-02-18" nation="" />
     <ATHLETE firstname="Ari-Pekka" nameprefix="" lastname="Liukkonen" gender="M" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:00:48.72">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-05-26" nation="" />
     <ATHLETE firstname="Vladislav" nameprefix="" lastname="Grinev" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:50.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-16" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Durango" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:04:00.96">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-06-05" nation="" />
     <ATHLETE firstname="Alexander" nameprefix="" lastname="Fedorov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:08:24.46">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-12" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Heron" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:15:49.04">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-12" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Heron" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:25.44">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2016-04-03" nation="" />
     <ATHLETE firstname="Anton" nameprefix="" lastname="Butymov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:55.09">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-11-21" nation="" />
     <ATHLETE firstname="Ryota" nameprefix="" lastname="Maejima" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:02.76">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-04-26" nation="" />
     <ATHLETE firstname="Dmitri" nameprefix="" lastname="Gorbunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:27.21">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-04-18" nation="" />
     <ATHLETE firstname="Kirill" nameprefix="" lastname="Strelnikov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:00.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-04-16" nation="" />
     <ATHLETE firstname="Kirill" nameprefix="" lastname="Strelnikov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:11.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2013-08-10" nation="" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Burckle" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:23.71">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2008-08-16" nation="" />
     <ATHLETE firstname="Kohei" nameprefix="" lastname="Kawamoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:53.09">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2008-08-15" nation="" />
     <ATHLETE firstname="Kohei" nameprefix="" lastname="Kawamoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:00.74">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-06-05" nation="" />
     <ATHLETE firstname="Aleksandr" nameprefix="" lastname="Pribytok" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:03.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-04-28" nation="" />
     <ATHLETE firstname="Dmitri" nameprefix="" lastname="Gorbunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:04:30.05">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-09-12" nation="" />
     <ATHLETE firstname="Diogo" nameprefix="" lastname="Yabe" gender="M" nation="BRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:23.49">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Blue Marlins (SG)" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:00:52.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Blue Marlins (SG)" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:01:58.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-09-03" nation="NED" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Oosting" gender="M" nation="NED" CLUB="PSV" birthdate="1981-04-01" />
    </RECORD>
    <RECORD swimtime="00:04:14.13">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Londen" date="2016-05-25" nation="GBR" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:08:41.84">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Londen" date="2016-05-25" nation="GBR" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:17:17.26">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2015-05-08" nation="NED" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Schr�der" gender="M" nation="NED" CLUB="TriVia" birthdate="1984-09-16" />
    </RECORD>
    <RECORD swimtime="00:00:27.89">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2017-05-05" nation="NED" />
     <ATHLETE firstname="Dirk" nameprefix="" lastname="Gielink" gender="M" nation="NED" CLUB="Aqua-Novio&apos;94" birthdate="1983-02-03" />
    </RECORD>
    <RECORD swimtime="00:01:03.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <ATHLETE firstname="Joan" nameprefix="" lastname="Kentrop" gender="M" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1985-12-01" />
    </RECORD>
    <RECORD swimtime="00:02:18.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2012-05-04" nation="NED" />
     <ATHLETE firstname="Dennis" nameprefix="" lastname="Brouwers" gender="M" nation="NED" CLUB="HZPC" birthdate="1978-07-14" />
    </RECORD>
    <RECORD swimtime="00:00:30.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Joan" nameprefix="" lastname="Kentrop" gender="M" nation="NED" CLUB="Aquarijn" birthdate="1985-12-01" />
    </RECORD>
    <RECORD swimtime="00:01:07.12">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2011-05-08" nation="NED" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Claus" gender="M" nation="NED" CLUB="Heldense Zwemvereniging" birthdate="1980-04-28" />
    </RECORD>
    <RECORD swimtime="00:02:32.94">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Den Haag" date="2014-05-03" nation="NED" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Claus" gender="M" nation="NED" CLUB="Swimteam Helden-Mosa" birthdate="1980-04-28" />
    </RECORD>
    <RECORD swimtime="00:00:25.32">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Blue Marlins (SG)" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:00:56.58">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" CLUB="Blue Marlins (SG)" birthdate="1992-08-21" />
    </RECORD>
    <RECORD swimtime="00:02:17.79">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Matteo" nameprefix="" lastname="Viani" gender="M" nation="NED" CLUB="Zwemlust-den Hommel" birthdate="1990-06-22" />
    </RECORD>
    <RECORD swimtime="00:02:15.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Prague" date="1997-09-07" nation="CZE" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:57.25">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Apeldoorn" date="1995-06-10" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:22.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Jyv�skyl�" date="2020-02-15" nation="FIN" />
     <ATHLETE firstname="Ari-Pekka" nameprefix="" lastname="Liukkonen" gender="M" nation="FIN" />
    </RECORD>
    <RECORD swimtime="00:00:50.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="St. Petersburg" date="2018-06-03" nation="RUS" />
     <ATHLETE firstname="Evgeni" nameprefix="" lastname="Lagunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:53.33">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="G�teborg" date="2010-08-02" nation="SWE" />
     <ATHLETE firstname="Jacob" nameprefix="" lastname="Carstensen" gender="M" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:04:01.70">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2012-06-16" nation="ITA" />
     <ATHLETE firstname="Jacob" nameprefix="" lastname="Carstensen" gender="M" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:08:08.53">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-11" nation="GER" />
     <ATHLETE firstname="Jan" nameprefix="" lastname="Wolfgarten" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:15:25.79">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-11" nation="GER" />
     <ATHLETE firstname="Jan" nameprefix="" lastname="Wolfgarten" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:26.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Leipzig" date="2011-05-07" nation="GER" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Herbst" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:56.55">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Leipzig" date="2011-05-07" nation="GER" />
     <ATHLETE firstname="Stefan" nameprefix="" lastname="Herbst" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:04.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="G�teborg" date="2010-08-01" nation="SWE" />
     <ATHLETE firstname="Razvan" nameprefix="" lastname="Florea" gender="M" nation="ROU" />
    </RECORD>
    <RECORD swimtime="00:00:28.24">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kazan" date="2015-08-13" nation="RUS" />
     <ATHLETE firstname="Sergei" nameprefix="" lastname="Geibel" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:03.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="London" date="2016-05-27" nation="GBR" />
     <ATHLETE firstname="Wolfgang" nameprefix="" lastname="Maier" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:18.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2022-04-23" nation="RUS" />
     <ATHLETE firstname="Dmitri" nameprefix="" lastname="Gorbunov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:24.25">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Obninsk" date="2018-04-28" nation="RUS" />
     <ATHLETE firstname="Nikita" nameprefix="" lastname="Konovalov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:54.12">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-17" nation="HUN" />
     <ATHLETE firstname="Maxim" nameprefix="" lastname="Ganikhin" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:05.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Maxim" nameprefix="" lastname="Ganikhin" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:07.38">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="G�teborg" date="2010-08-03" nation="SWE" />
     <ATHLETE firstname="Jacob" nameprefix="" lastname="Carstensen" gender="M" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:04:24.11">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="W�rzburg" date="2013-03-09" nation="GER" />
     <ATHLETE firstname="Lukasz" nameprefix="" lastname="Wojt" gender="M" nation="POL" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="30" agemax="34" />
   <RECORDS>
    <RECORD swimtime="00:00:22.13">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2013-07-13" nation="" />
     <ATHLETE firstname="Roland" nameprefix="" lastname="Schoeman" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:49.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-07-23" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:49.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-08-06" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:58.12">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-07-23" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:08.53">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-11" nation="GER" />
     <ATHLETE firstname="Jan" nameprefix="" lastname="Wolfgarten" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:15:25.79">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-11" nation="GER" />
     <ATHLETE firstname="Jan" nameprefix="" lastname="Wolfgarten" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:25.53">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-09-24" nation="" />
     <ATHLETE firstname="Sergey" nameprefix="" lastname="Fesikov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:55.93">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2014-07-13" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:02.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2000-11-24" nation="" />
     <ATHLETE firstname="Rogerio" nameprefix="" lastname="Romero" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:00:27.74">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-03-12" nation="" />
     <ATHLETE firstname="Kohhei" nameprefix="" lastname="Tominaga" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:01.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-08-31" nation="" />
     <ATHLETE firstname="Ryo" nameprefix="" lastname="Kobayashi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:16.79">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-08-10" nation="" />
     <ATHLETE firstname="Shotaro" nameprefix="" lastname="Shimazaki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:23.16">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-05-26" nation="" />
     <ATHLETE firstname="Oleg" nameprefix="" lastname="Kostin" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:53.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-04-08" nation="" />
     <ATHLETE firstname="Henrique" nameprefix="" lastname="Martins" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:02:03.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-08-17" nation="" />
     <ATHLETE firstname="Takatsugu" nameprefix="" lastname="Oga" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:02.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-05-22" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:20.81">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-07-23" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:24.76">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Londen" date="2016-05-29" nation="GBR" />
     <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" CLUB="d&apos;ELFT" birthdate="1980-05-09" />
    </RECORD>
    <RECORD swimtime="00:00:53.87">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Londen" date="2016-05-28" nation="GBR" />
     <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" CLUB="d&apos;ELFT" birthdate="1980-05-09" />
    </RECORD>
    <RECORD swimtime="00:01:59.61">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Munchen" date="2000-08-02" nation="GER" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC " birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:20.44">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Innsbruck" date="1999-08-29" nation="AUT" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:09:11.35">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Remco" nameprefix="van" lastname="Althuis" gender="M" nation="NED" CLUB="PSV" birthdate="1983-01-25" />
    </RECORD>
    <RECORD swimtime="00:17:39.55">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-03" nation="NED" />
     <ATHLETE firstname="Remco" nameprefix="van" lastname="Althuis" gender="M" nation="NED" CLUB="PSV" birthdate="1983-01-25" />
    </RECORD>
    <RECORD swimtime="00:00:28.83">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2007-04-21" nation="NED" />
     <ATHLETE firstname="Theo Jan" nameprefix="" lastname="Tanis" gender="M" nation="NED" CLUB="De Gooye" birthdate="1969-03-16" />
    </RECORD>
    <RECORD swimtime="00:01:03.01">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1980-05-09" />
    </RECORD>
    <RECORD swimtime="00:02:16.14">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Londen" date="2016-05-28" nation="GBR" />
     <ATHLETE firstname="Dennis" nameprefix="" lastname="Brouwers" gender="M" nation="NED" CLUB="HZPC" birthdate="1978-07-14" />
    </RECORD>
    <RECORD swimtime="00:00:30.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-09-03" nation="NED" />
     <ATHLETE firstname="Martin" nameprefix="de" lastname="Wildt" gender="M" nation="NED" CLUB="Nuenen" birthdate="1974-03-16" />
    </RECORD>
    <RECORD swimtime="00:01:06.33">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Claus" gender="M" nation="NED" CLUB="Swimteam Helden-Mosa (SG)" birthdate="1980-04-28" />
    </RECORD>
    <RECORD swimtime="00:02:26.21">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-09-06" nation="NED" />
     <ATHLETE firstname="Martin" nameprefix="de" lastname="Wildt" gender="M" nation="NED" CLUB="Nuenen" birthdate="1974-03-16" />
    </RECORD>
    <RECORD swimtime="00:00:26.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Kampen" date="1999-04-17" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:59.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Palma de Mallorca" date="2001-07-04" nation="ESP" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:19.11">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="1996-06-27" nation="GBR" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:13.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Palma de Mallorca" date="2001-07-03" nation="ESP" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:54.18">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Munchen" date="2000-07-31" nation="GER" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC " birthdate="1963-04-24" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:22.76">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Stockholm" date="2005-08-20" nation="SWE" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Foster" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:51.52">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Reus" date="2018-07-07" nation="ESP" />
     <ATHLETE firstname="Mikel" nameprefix="" lastname="Bildosola Agirregomezkorta" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:55.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kazan" date="2015-08-12" nation="RUS" />
     <ATHLETE firstname="Ioan" nameprefix="" lastname="Gherghel" gender="M" nation="ROU" />
    </RECORD>
    <RECORD swimtime="00:04:05.91">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-10" nation="GER" />
     <ATHLETE firstname="Petar" nameprefix="" lastname="Stoychev" gender="M" nation="BUL" />
    </RECORD>
    <RECORD swimtime="00:08:18.44">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-12" nation="GER" />
     <ATHLETE firstname="Petar" nameprefix="" lastname="Stoychev" gender="M" nation="BUL" />
    </RECORD>
    <RECORD swimtime="00:16:00.04">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="W�rzburg" date="2012-03-11" nation="GER" />
     <ATHLETE firstname="Petar" nameprefix="" lastname="Stoychev" gender="M" nation="BUL" />
    </RECORD>
    <RECORD swimtime="00:00:26.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="London" date="2016-05-29" nation="GBR" />
     <ATHLETE firstname="Lubos" nameprefix="" lastname="Krizko" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:00:58.48">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Riccione" date="2016-06-25" nation="ITA" />
     <ATHLETE firstname="Marco" nameprefix="" lastname="Maccianti" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:07.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Riccione" date="2016-06-22" nation="ITA" />
     <ATHLETE firstname="Marco" nameprefix="" lastname="Maccianti" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:28.68">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kranj" date="2018-09-03" nation="SLO" />
     <ATHLETE firstname="Markic" nameprefix="" lastname="Matjaz" gender="M" nation="SLO" />
    </RECORD>
    <RECORD swimtime="00:01:02.72">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Vantaa" date="2009-10-25" nation="FIN" />
     <ATHLETE firstname="Vladislav" nameprefix="" lastname="Bragin" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:20.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Riccione" date="2004-06-05" nation="ITA" />
     <ATHLETE firstname="Nick" nameprefix="" lastname="Gillingham" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:24.38">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Magdeburg" date="2022-05-07" nation="GER" />
     <ATHLETE firstname="Stefano" nameprefix="" lastname="Razeto" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:54.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Obninsk" date="2019-04-28" nation="RUS" />
     <ATHLETE firstname="Nikolay" nameprefix="" lastname="Skvortsov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:02.54">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Obninsk" date="2019-04-26" nation="RUS" />
     <ATHLETE firstname="Nikolay" nameprefix="" lastname="Skvortsov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:09.85">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gwangju" date="2019-08-15" nation="KOR" />
     <ATHLETE firstname="Ioannis" nameprefix="" lastname="Drymonakos" gender="M" nation="GRE" />
    </RECORD>
    <RECORD swimtime="00:04:36.66">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gwangju" date="2019-08-14" nation="KOR" />
     <ATHLETE firstname="Ioannis" nameprefix="" lastname="Drymonakos" gender="M" nation="GRE" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="35" agemax="39" />
   <RECORDS>
    <RECORD swimtime="00:00:22.76">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Stockholm" date="2005-08-20" nation="SWE" />
     <ATHLETE firstname="Mark" nameprefix="" lastname="Foster" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:50.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-09-27" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Hara" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:51.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-07" nation="" />
     <ATHLETE firstname="Shogo" nameprefix="" lastname="Hirara" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:04:05.91">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2012-03-10" nation="" />
     <ATHLETE firstname="Petar" nameprefix="" lastname="Stoychev" gender="M" nation="BUL" />
    </RECORD>
    <RECORD swimtime="00:08:18.44">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2012-03-10" nation="" />
     <ATHLETE firstname="Petar" nameprefix="" lastname="Stoychev" gender="M" nation="BUL" />
    </RECORD>
    <RECORD swimtime="00:16:00.04">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2012-03-11" nation="" />
     <ATHLETE firstname="Petar" nameprefix="" lastname="Stoychev" gender="M" nation="BUL" />
    </RECORD>
    <RECORD swimtime="00:00:26.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-05-07" nation="" />
     <ATHLETE firstname="Stefano" nameprefix="" lastname="Razeto" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:57.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-10-22" nation="" />
     <ATHLETE firstname="Manabu" nameprefix="" lastname="Sasaki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:07.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2016-06-22" nation="" />
     <ATHLETE firstname="Marco" nameprefix="" lastname="Maccianti" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.83">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-08-11" nation="" />
     <ATHLETE firstname="Ryouta" nameprefix="" lastname="Nomura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:02.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2020-02-11" nation="JPN" />
     <ATHLETE firstname="Ryo" nameprefix="" lastname="Kobayashi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:20.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Riccione" date="2004-06-05" nation="ITA" />
     <ATHLETE firstname="Nick" nameprefix="" lastname="Gillingham" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:24.03">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-12-02" nation="" />
     <ATHLETE firstname="Benjamin" nameprefix="" lastname="Hockin" gender="M" nation="PAR" />
    </RECORD>
    <RECORD swimtime="00:00:53.65">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2018-08-02" nation="" />
     <ATHLETE firstname="Kohei" nameprefix="" lastname="Kawamoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:02.54">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2019-04-26" nation="" />
     <ATHLETE firstname="Nikolay" nameprefix="" lastname="Skvortsov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:05.65">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-07-07" nation="" />
     <ATHLETE firstname="Darian" nameprefix="" lastname="Townsend" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:36.66">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-08-14" nation="" />
     <ATHLETE firstname="Ioannis" nameprefix="" lastname="Drymonakos" gender="M" nation="GRE" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:24.76">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:00:54.42">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:02:02.01">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Millau" date="2003-08-27" nation="FRA" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:04:28.16">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Stockholm" date="2005-08-19" nation="SWE" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:09:21.92">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Cadiz" date="2009-09-15" nation="ESP" />
     <ATHLETE firstname="Joost" nameprefix="" lastname="Kuijlaars" gender="M" nation="NED" CLUB="MNC Dordrecht" birthdate="1966-01-01" />
    </RECORD>
    <RECORD swimtime="00:17:46.39">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Apeldoorn" date="2006-06-11" nation="NED" />
     <ATHLETE firstname="Joost" nameprefix="" lastname="Kuijlaars" gender="M" nation="NED" CLUB="MNC Dordrecht" birthdate="1966-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:28.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2009-05-10" nation="NED" />
     <ATHLETE firstname="Theo Jan" nameprefix="" lastname="Tanis" gender="M" nation="NED" CLUB="De Schotejil" birthdate="1969-03-16" />
    </RECORD>
    <RECORD swimtime="00:01:03.21">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2011-05-07" nation="NED" />
     <ATHLETE firstname="Theo Jan" nameprefix="" lastname="Tanis" gender="M" nation="NED" CLUB="De Schotejil" birthdate="1969-03-16" />
    </RECORD>
    <RECORD swimtime="00:02:19.85">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Dennis" nameprefix="" lastname="Brouwers" gender="M" nation="NED" CLUB="HZPC" birthdate="1978-07-14" />
    </RECORD>
    <RECORD swimtime="00:00:30.77">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Luxembourg" date="2009-10-17" nation="LUX" />
     <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" CLUB="PSV" birthdate="1968-10-13" />
    </RECORD>
    <RECORD swimtime="00:01:07.54">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kranj" date="2018-09-07" nation="SLO" />
     <ATHLETE firstname="Martin" nameprefix="de" lastname="Wildt" gender="M" nation="NED" CLUB="Nuenen" birthdate="1974-03-16" />
    </RECORD>
    <RECORD swimtime="00:02:28.07">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Martin" nameprefix="de" lastname="Wildt" gender="M" nation="NED" CLUB="Nuenen" birthdate="1974-03-16" />
    </RECORD>
    <RECORD swimtime="00:00:26.66">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Apeldoorn" date="2003-06-15" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:01:00.82">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Luxembourg" date="2003-10-18" nation="LUX" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:18.45">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Portland" date="1998-08-11" nation="USA" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:19.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Millau" date="2003-08-26" nation="FRA" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:05:00.37">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2016-05-07" nation="NED" />
     <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" CLUB="d&apos;ELFT WAVE (SG)" birthdate="1976-06-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:23.14">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Barcelona" date="2023-06-03" nation="ESP" />
     <ATHLETE firstname="Mikel" nameprefix="" lastname="Bildosola Agirregomezkorta" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:50.73">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2023-06-30" nation="ITA" />
     <ATHLETE firstname="Filipo" nameprefix="" lastname="Magnini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:55.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-16" nation="HUN" />
     <ATHLETE firstname="Claus" nameprefix="" lastname="Iversen" gender="M" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:04:08.67">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gwangju" date="2019-08-18" nation="KOR" />
     <ATHLETE firstname="Nicola" nameprefix="" lastname="Nisato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:08:35.85">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gwangju" date="2019-08-12" nation="KOR" />
     <ATHLETE firstname="Nicola" nameprefix="" lastname="Nisato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:16:24.76">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Lodi" date="2018-04-07" nation="ITA" />
     <ATHLETE firstname="Nicola" nameprefix="" lastname="Nisato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Genova" date="2009-02-01" nation="ITA" />
     <ATHLETE firstname="Giuseppe" nameprefix="" lastname="Tiano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:59.24">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Riccione" date="2023-07-01" nation="ITA" />
     <ATHLETE firstname="Enrico" nameprefix="" lastname="Catalano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:10.46">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="London" date="2016-05-28" nation="GBR" />
     <ATHLETE firstname="Maurizio" nameprefix="" lastname="Tersar" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:28.84">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Cadiz" date="2009-09-16" nation="ESP" />
     <ATHLETE firstname="Alberto" nameprefix="" lastname="Montini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:03.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2012-05-20" nation="RUS" />
     <ATHLETE firstname="Vladislav" nameprefix="" lastname="Bragin" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:22.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Riccione " date="2012-06-15" nation="ITA" />
     <ATHLETE firstname="Alberto" nameprefix="" lastname="Montini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:24.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-07" nation="JPN" />
     <ATHLETE firstname="Andrejs" nameprefix="" lastname="Duda" gender="M" nation="LAT" />
    </RECORD>
    <RECORD swimtime="00:00:55.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-08" nation="JPN" />
     <ATHLETE firstname="Andrejs" nameprefix="" lastname="Duda" gender="M" nation="LAT" />
    </RECORD>
    <RECORD swimtime="00:02:09.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Claus" nameprefix="" lastname="Iversen" gender="M" nation="DEN" />
    </RECORD>
    <RECORD swimtime="00:02:11.67">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Cadiz" date="2009-09-15" nation="ESP" />
     <ATHLETE firstname="Alberto" nameprefix="" lastname="Montini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:04:43.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Riccione" date="2012-06-12" nation="ITA" />
     <ATHLETE firstname="Uwe" nameprefix="" lastname="Volk" gender="M" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="40" agemax="44" />
   <RECORDS>
    <RECORD swimtime="00:00:23.14">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-08" nation="" />
     <ATHLETE firstname="Andrei" nameprefix="" lastname="Kurnosov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:50.73">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-06-30" nation="" />
     <ATHLETE firstname="Filippo" nameprefix="" lastname="Magnini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:53.65">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2010-08-02" nation="" />
     <ATHLETE firstname="Vladimir" nameprefix="" lastname="Pyshnenko" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:06.74">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-07-24" nation="" />
     <ATHLETE firstname="Erik" nameprefix="" lastname="Hochstein" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:35.85">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-12-08" nation="" />
     <ATHLETE firstname="Nicola" nameprefix="" lastname="Nisato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:16:24.76">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-04-07" nation="" />
     <ATHLETE firstname="Nicola" nameprefix="" lastname="Nisato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.13">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-08-18" nation="" />
     <ATHLETE firstname="Nicholas" nameprefix="" lastname="Neckles" gender="M" nation="BAR" />
    </RECORD>
    <RECORD swimtime="00:00:58.45">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-08-17" nation="" />
     <ATHLETE firstname="Nicholas" nameprefix="" lastname="Neckles" gender="M" nation="BAR" />
    </RECORD>
    <RECORD swimtime="00:02:08.06">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-08-13" nation="" />
     <ATHLETE firstname="Nicholas" nameprefix="" lastname="Neckles" gender="M" nation="BAR" />
    </RECORD>
    <RECORD swimtime="00:00:28.84">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Cadiz" date="2009-09-16" nation="ESP" />
     <ATHLETE firstname="Alberto" nameprefix="" lastname="Montini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:03.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2012-05-20" nation="RUS" />
     <ATHLETE firstname="Vladislav" nameprefix="" lastname="Bragin" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:18.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2015-07-11" nation="" />
     <ATHLETE firstname="Steven" nameprefix="" lastname="West" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:24.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-07" nation="" />
     <ATHLETE firstname="Andrejs" nameprefix="" lastname="Duda" gender="M" nation="LAT" />
    </RECORD>
    <RECORD swimtime="00:00:55.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-05-20" nation="" />
     <ATHLETE firstname="Carlos" nameprefix="" lastname="Nascimento" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:02:05.55">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2004-07-11" nation="" />
     <ATHLETE firstname="Dennis" nameprefix="" lastname="Baker" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:08.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-05-27" nation="" />
     <ATHLETE firstname="Markus" nameprefix="" lastname="Rogan" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:43.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Riccione" date="2012-06-12" nation="ITA" />
     <ATHLETE firstname="Uwe" nameprefix="" lastname="Volk" gender="M" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:25.22">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2009-03-22" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:55.69">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:02:05.03">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:04:35.06">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2009-03-22" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:09:46.04">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg" date="2018-10-14" nation="LUX" />
     <ATHLETE firstname="Pieter" nameprefix="van" lastname="Gemeren" gender="M" nation="NED" CLUB="DAW" birthdate="1969-10-21" />
    </RECORD>
    <RECORD swimtime="00:18:59.27">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg" date="2018-10-13" nation="LUX" />
     <ATHLETE firstname="Pieter" nameprefix="van" lastname="Gemeren" gender="M" nation="NED" CLUB="DAW" birthdate="1969-10-21" />
    </RECORD>
    <RECORD swimtime="00:00:29.36">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2009-03-22" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:01:05.82">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Tjakko" nameprefix="" lastname="Ruinemans" gender="M" nation="NED" CLUB="De Dinkel" birthdate="1974-08-23" />
    </RECORD>
    <RECORD swimtime="00:02:20.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Cadiz" date="2009-09-18" nation="ESP" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:31.82">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Joost" nameprefix="" lastname="Hoetjes" gender="M" nation="NED" CLUB="DAW" birthdate="1978-07-19" />
    </RECORD>
    <RECORD swimtime="00:01:10.52">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Joost" nameprefix="" lastname="Hoetjes" gender="M" nation="NED" CLUB="DAW" birthdate="1978-07-19" />
    </RECORD>
    <RECORD swimtime="00:02:37.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Cadiz" date="2009-09-19" nation="ESP" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:27.09">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1978-10-02" />
    </RECORD>
    <RECORD swimtime="00:01:00.64">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Cadiz" date="2009-09-16" nation="ESP" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:17.94">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2007-04-21" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:18.80">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Cadiz" date="2009-09-15" nation="ESP" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:05:07.68">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2008-01-18" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:23.98">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Olympic" date="2014-07-05" nation="RUS" />
     <ATHLETE firstname="Vladimir" nameprefix="" lastname="Predkin" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:53.66">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-15" nation="HUN" />
     <ATHLETE firstname="Valter" nameprefix="" lastname="Kalaus" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:01:57.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Montreal" date="2014-08-05" nation="CAN" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:13.86">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2012-06-16" nation="ITA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:08:40.79">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kazan" date="2015-08-10" nation="RUS" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:16:42.01">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Lignano" date="2023-02-03" nation="ITA" />
     <ATHLETE firstname="Nicola" nameprefix="" lastname="Nisato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.62">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="St. Petersburg" date="2021-06-05" nation="RUS" />
     <ATHLETE firstname="Alexandr" nameprefix="" lastname="Shilin" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:00.97">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Serkan" nameprefix="" lastname="Atasay" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:02:13.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Riccione" date="2023-06-28" nation="ITA" />
     <ATHLETE firstname="Maurizio" nameprefix="" lastname="Tersar" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:29.51">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-20" nation="HUN" />
     <ATHLETE firstname="Serkan" nameprefix="" lastname="Atasay" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:01:05.33">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="London" date="2016-05-27" nation="GBR" />
     <ATHLETE firstname="Vladislav" nameprefix="" lastname="Bragin" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:24.39">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Treviso" date="2013-05-31" nation="ITA" />
     <ATHLETE firstname="Alberto" nameprefix="" lastname="Montini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:25.48">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-16" nation="HUN" />
     <ATHLETE firstname="Serkan" nameprefix="" lastname="Atasay" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:00:57.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Budapest" date="2017-08-17" nation="HUN" />
     <ATHLETE firstname="Serkan" nameprefix="" lastname="Atasay" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:02:13.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Legnano" date="2019-02-02" nation="ITA" />
     <ATHLETE firstname="Andrea" nameprefix="" lastname="Marcato" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:10.24">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Zaragoza" date="2015-07-25" nation="ESP" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:43.83">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Montreal " date="2014-08-05" nation="CAN" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="45" agemax="49" />
   <RECORDS>
    <RECORD swimtime="00:00:23.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-08-15" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Hara" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:52.24">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-08-13" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Hara" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:57.75">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Montreal" date="2014-08-05" nation="CAN" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:11.07">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-08-09" nation="" />
     <ATHLETE firstname="Keith" nameprefix="" lastname="Switzer" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:40.79">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-08-10" nation="" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:16:38.81">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-08-10" nation="" />
     <ATHLETE firstname="Jeff" nameprefix="" lastname="Erwin" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:27.56">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-06-04" nation="" />
     <ATHLETE firstname="Marcin" nameprefix="" lastname="Kaczmarek" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:00:59.57">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-08-04" nation="" />
     <ATHLETE firstname="Chuck" nameprefix="" lastname="Barnes" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:11.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2013-06-07" nation="" />
     <ATHLETE firstname="Eduardo" nameprefix="" lastname="Marocco" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:00:29.22">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-08-09" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Togo" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:04.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-07-14" nation="" />
     <ATHLETE firstname="Steven" nameprefix="" lastname="West" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:19.44">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2018-06-22" nation="" />
     <ATHLETE firstname="Steven" nameprefix="" lastname="West" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:25.07">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-07" nation="" />
     <ATHLETE firstname="Marc Kevin" nameprefix="" lastname="Allan" gender="M" nation="RSA" />
    </RECORD>
    <RECORD swimtime="00:00:56.85">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2002-08-11" nation="" />
     <ATHLETE firstname="Paul" nameprefix="" lastname="Carter" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:06.94">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2006-08-09" nation="" />
     <ATHLETE firstname="Dennis" nameprefix="" lastname="Baker" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:10.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-08-07" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:43.83">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2014-08-05" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:26.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:00:57.05">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-09-05" nation="NED" />
     <ATHLETE firstname="Cees" nameprefix="van" lastname="Houwelingen" gender="M" nation="NED" CLUB="De Schelde" birthdate="1963-03-24" />
    </RECORD>
    <RECORD swimtime="00:02:08.84">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-05-10" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:04:40.35">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Dordrecht" date="2012-04-01" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:09:46.85">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Casablanca" date="1998-06-25" nation="MAR" />
     <ATHLETE firstname="Donald" nameprefix="" lastname="Uijtenbogaart" gender="M" nation="NED" CLUB="De Dolfijn" birthdate="1947-01-01" />
    </RECORD>
    <RECORD swimtime="00:18:50.20">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-02" nation="NED" />
     <ATHLETE firstname="Bob" nameprefix="de" lastname="Vries" gender="M" nation="NED" CLUB="The Hague Swimming (SG)" birthdate="1966-04-13" />
    </RECORD>
    <RECORD swimtime="00:00:29.78">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1969-11-26" />
    </RECORD>
    <RECORD swimtime="00:01:06.23">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2014-05-03" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:25.16">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Londen" date="2016-05-28" nation="GBR" />
     <ATHLETE firstname="Jan Gert" nameprefix="" lastname="Notenbomer" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1966-08-04" />
    </RECORD>
    <RECORD swimtime="00:00:32.96">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" CLUB="PSV" birthdate="1968-10-13" />
    </RECORD>
    <RECORD swimtime="00:01:13.93">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Alkmaar" date="2017-04-09" nation="NED" />
     <ATHLETE firstname="Jan Gert" nameprefix="" lastname="Notenbomer" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1966-08-04" />
    </RECORD>
    <RECORD swimtime="00:02:42.82">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-09-06" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:00:27.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2009-05-10" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:00:59.67">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2009-05-10" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:15.06">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2009-05-09" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:24.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2013-09-02" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="AZ&amp;PC" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:05:06.60">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2009-05-08" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:24.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Obninsk" date="2019-04-27" nation="RUS" />
     <ATHLETE firstname="Vladimir" nameprefix="" lastname="Predkin" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:54.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vichy" date="2017-06-30" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:58.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vichy" date="2017-07-01" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:17.28">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Vichy" date="2017-06-30" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:08:49.22">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kranj" date="2018-09-02" nation="SLO" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:17:35.40">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Napoli" date="2018-06-10" nation="ITA" />
     <ATHLETE firstname="Dino" nameprefix="" lastname="Schorn" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:28.64">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Vichy" date="2017-06-30" nation="FRA" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:03.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Roma" date="2022-09-02" nation="ITA" />
     <ATHLETE firstname="Frank" nameprefix="" lastname="Gruner" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:16.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Fukuoka" date="2023-08-06" nation="JPN" />
     <ATHLETE firstname="Frank" nameprefix="" lastname="Gruner" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:30.16">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2021-06-05" nation="RUS" />
     <ATHLETE firstname="Vladislav" nameprefix="" lastname="Bragin" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:06.14">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2022-04-22" nation="RUS" />
     <ATHLETE firstname="Vladislav" nameprefix="" lastname="Bragin" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:02:25.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2022-04-23" nation="RUS" />
     <ATHLETE firstname="Vladislav" nameprefix="" lastname="Bragin" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:00:25.98">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Coque" date="2023-07-08" nation="LUX" />
     <ATHLETE firstname="Fr�d�ric" nameprefix="" lastname="Tonus" gender="M" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:00:58.62">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Fr�d�ric" nameprefix="" lastname="Tonus" gender="M" nation="BEL" />
    </RECORD>
    <RECORD swimtime="00:02:14.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Kazan" date="2015-08-15" nation="RUS" />
     <ATHLETE firstname="Mauro" nameprefix="" lastname="Cappelletti" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:13.96">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Kranj" date="2018-09-05" nation="SLO" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:50.33">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Charleroi" date="2017-04-15" nation="BEL" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="50" agemax="54" />
   <RECORDS>
    <RECORD swimtime="00:00:24.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-06-27" nation="" />
     <ATHLETE firstname="Brent" nameprefix="" lastname="Barnes" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:54.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-06-30" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:58.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-01-07" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:15.93">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-04" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:08:55.05">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2010-07-31" nation="" />
     <ATHLETE firstname="Marcus" nameprefix="" lastname="Mattioli" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:17:08.33">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2000-08-20" nation="" />
     <ATHLETE firstname="Jim" nameprefix="" lastname="McConica" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.20">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-05-28" nation="" />
     <ATHLETE firstname="M." nameprefix="" lastname="Gromov-Ivanov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:01.57">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-08-06" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:02:14.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-08-05" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:29.70">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-08-11" nation="" />
     <ATHLETE firstname="Hideaki" nameprefix="" lastname="Togo" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:06.12">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-07-10" nation="" />
     <ATHLETE firstname="Steve" nameprefix="" lastname="West" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:24.44">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-07-09" nation="" />
     <ATHLETE firstname="Steve" nameprefix="" lastname="West" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:25.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-05-20" nation="" />
     <ATHLETE firstname="Serkan" nameprefix="" lastname="Atasay" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:00:56.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-08" nation="" />
     <ATHLETE firstname="Eiji" nameprefix="" lastname="Nomura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:13.26">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-11-06" nation="" />
     <ATHLETE firstname="Eiji" nameprefix="" lastname="Nomura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:11.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-08-06" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:04:45.61">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-08-03" nation="" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:26.43">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:00:59.55">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-05-04" nation="NED" />
     <ATHLETE firstname="Albert" nameprefix="" lastname="Boonstra" gender="M" nation="NED" CLUB="Aqua-Novio&apos;94" birthdate="1957-05-22" />
    </RECORD>
    <RECORD swimtime="00:02:10.32">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-02" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:04:39.18">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-09-02" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:09:39.03">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-02" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:18:41.25">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-04" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:00:31.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Riccione" date="2012-06-16" nation="ITA" />
     <ATHLETE firstname="Albert" nameprefix="" lastname="Boonstra" gender="M" nation="NED" CLUB="Aqua-Novio&apos;94" birthdate="1957-05-22" />
    </RECORD>
    <RECORD swimtime="00:01:09.36">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:02:29.06">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2013-09-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:00:33.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Antwerpen" date="2023-02-05" nation="BEL" />
     <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" CLUB="PSV" birthdate="1968-10-13" />
    </RECORD>
    <RECORD swimtime="00:01:16.78">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Copenhagen" date="2009-07-29" nation="DEN" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:02:47.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="Jan Gert" nameprefix="" lastname="Notenbomer" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1966-08-04" />
    </RECORD>
    <RECORD swimtime="00:00:27.47">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2013-09-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:01.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2013-09-03" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:19.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2013-05-04" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:25.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2013-09-02" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:05:22.27">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2015-05-10" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="Albion" birthdate="1958-09-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:25.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Fukuoka" date="2023-08-09" nation="JPN" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Hodgson" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:56.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kranj" date="2018-09-06" nation="SLO" />
     <ATHLETE firstname="Ahmet" nameprefix="" lastname="Nakkas" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:02:04.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-16" nation="HUN" />
     <ATHLETE firstname="Ahmet" nameprefix="" lastname="Nakkas" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:04:31.94">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Fukuoka" date="2023-08-11" nation="JPN" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Dixon" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:09:12.59">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Fukuoka" date="2023-08-05" nation="JPN" />
     <ATHLETE firstname="Fabio" nameprefix="" lastname="Calmasini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:18:00.36">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Trevisio" date="2022-05-20" nation="ITA" />
     <ATHLETE firstname="Luca" nameprefix="di" lastname="Iacovo" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:30.15">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Hodgson" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:04.84">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Fukuoka" date="2023-08-10" nation="JPN" />
     <ATHLETE firstname="Alessio" nameprefix="" lastname="Germani" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:22.56">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Roma" date="2022-09-01" nation="ITA" />
     <ATHLETE firstname="Alessio" nameprefix="" lastname="Germani" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:30.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Torino" date="2019-06-02" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:07.65">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Gwangju" date="2019-08-13" nation="KOR" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:30.67">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Palermo" date="2018-07-11" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:26.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-07" nation="JPN" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Hodgson" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:01.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2013-09-03" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:19.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2013-05-04" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:19.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Rades" date="2023-05-10" nation="TUN" />
     <ATHLETE firstname="Nicolas" nameprefix="" lastname="Granger" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:05:14.38">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Roma" date="2022-08-30" nation="ITA" />
     <ATHLETE firstname="Antonella" nameprefix="" lastname="Laveglia" gender="M" nation="ITA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="55" agemax="59" />
   <RECORDS>
    <RECORD swimtime="00:00:24.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-07-19" nation="" />
     <ATHLETE firstname="Brent" nameprefix="" lastname="Barnes" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:56.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-02-24" nation="" />
     <ATHLETE firstname="Calvin" nameprefix="" lastname="Maughan" gender="M" nation="rsa" />
    </RECORD>
    <RECORD swimtime="00:02:04.01">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-07-26" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:22.49">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-07-25" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:00.09">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-07-24" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:22.61">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-08-10" nation="" />
     <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:29.03">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2016-08-20" nation="" />
     <ATHLETE firstname="Steve" nameprefix="" lastname="Wood" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:03.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2015-06-21" nation="" />
     <ATHLETE firstname="Steve" nameprefix="" lastname="Wood" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:20.83">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-07-20" nation="" />
     <ATHLETE firstname="Rip" nameprefix="" lastname="Esselstyn" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:30.02">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-02-06" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:07.65">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2019-08-13" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:30.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-08-21" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Guthrie" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:26.56">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-10-10" nation="" />
     <ATHLETE firstname="Steve" nameprefix="" lastname="Hiltabiddle" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:00.56">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2012-08-11" nation="" />
     <ATHLETE firstname="Paul" nameprefix="" lastname="Carter" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:16.78">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2015-08-15" nation="" />
     <ATHLETE firstname="Marcus" nameprefix="" lastname="Mattioli" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:02:20.67">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2020-02-22" nation="USA" />
     <ATHLETE firstname="Jerome" nameprefix="" lastname="Frentsos" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:57.55">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-04-02" nation="" />
     <ATHLETE firstname="Brent" nameprefix="" lastname="Foster" gender="M" nation="NZL" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:27.13">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:01:00.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:02:13.47">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:04:46.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Alkmaar" date="2018-04-08" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:10:03.69">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:19:08.78">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-02" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:00:32.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:01:10.93">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" CLUB="De Rog" birthdate="1963-02-23" />
    </RECORD>
    <RECORD swimtime="00:02:36.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Rome" date="2022-09-01" nation="ITA" />
     <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1962-02-13" />
    </RECORD>
    <RECORD swimtime="00:00:37.50">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Londen" date="2016-05-26" nation="GBR" />
     <ATHLETE firstname="Paul" nameprefix="" lastname="Bunnik" gender="M" nation="NED" CLUB="Triton" birthdate="1956-07-28" />
    </RECORD>
    <RECORD swimtime="00:01:21.89">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" CLUB="ZPC AMERSFOORT" birthdate="1963-04-24" />
    </RECORD>
    <RECORD swimtime="00:02:56.77">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2012-06-29" nation="HUN" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:00:27.65">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:02.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:23.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:31.35">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Kranj" date="2018-09-05" nation="SLO" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:05:31.07">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Gwangju" date="2019-08-14" nation="KOR" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="Albion d&apos;ELFT (SG)" birthdate="1958-09-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:26.00">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-17" nation="HUN" />
     <ATHLETE firstname="Alexey" nameprefix="" lastname="Markovskiy" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:57.66">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Roma" date="2022-09-04" nation="ITA" />
     <ATHLETE firstname="Ahmet" nameprefix="" lastname="Nakkas" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:02:08.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Las Palmas" date="2023-06-19" nation="ESP" />
     <ATHLETE firstname="Juan Carlos" nameprefix="" lastname="Vallejo Arroyo" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:04:30.15">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Las Palmas" date="2023-06-19" nation="ESP" />
     <ATHLETE firstname="Juan Carlos" nameprefix="" lastname="Vallejo Arroyo" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:09:39.23">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2016-06-21" nation="ITA" />
     <ATHLETE firstname="Marco" nameprefix="" lastname="Bravi" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:18:36.36">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Halle" date="2023-02-24" nation="GER" />
     <ATHLETE firstname="Karsten" nameprefix="" lastname="Dellbr�gge" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:31.18">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Aberdeen" date="2022-06-18" nation="GBR" />
     <ATHLETE firstname="Alec" nameprefix="" lastname="Johnson" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:07.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="St. Petersburg" date="2017-06-03" nation="RUS" />
     <ATHLETE firstname="Vladimir" nameprefix="" lastname="Gorkov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:29.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Obninsk" date="2018-04-27" nation="RUS" />
     <ATHLETE firstname="Vladimir" nameprefix="" lastname="Gorkov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:30.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Riccione" date="2023-06-30" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:09.57">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Fukuoka" date="2023-08-06" nation="JPN" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:33.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Riccione" date="2023-06-29" nation="ITA" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Sheffield" date="2023-06-04" nation="GBR" />
     <ATHLETE firstname="David" nameprefix="" lastname="Emerson" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:02.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:23.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:24.91">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Fukuoka" date="2023-08-08" nation="JPN" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:05:29.55">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Riccione" date="2012-06-12" nation="ITA" />
     <ATHLETE firstname="Lorenzo" nameprefix="" lastname="Marugo" gender="M" nation="ITA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="60" agemax="64" />
   <RECORDS>
    <RECORD swimtime="00:00:25.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2006-08-07" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:57.66">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-09-04" nation="" />
     <ATHLETE firstname="Ahmet" nameprefix="" lastname="Nakkas" gender="M" nation="TUR" />
    </RECORD>
    <RECORD swimtime="00:02:07.68">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-06" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Stephenson" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:30.15">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-06-19" nation="" />
     <ATHLETE firstname="Juan Carlos" nameprefix="" lastname="Vallejo Arroyo" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:09:21.08">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-05-20" nation="" />
     <ATHLETE firstname="Arnaldo" nameprefix="" lastname="Perez" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:55.91">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-03" nation="" />
     <ATHLETE firstname="Arnaldo" nameprefix="" lastname="Perez" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:30.59">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-10-08" nation="" />
     <ATHLETE firstname="Jamie" nameprefix="" lastname="Fowler" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:06.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-11-08" nation="" />
     <ATHLETE firstname="Jamie" nameprefix="" lastname="Fowler" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:26.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-08-08" nation="" />
     <ATHLETE firstname="Jamie" nameprefix="" lastname="Fowler" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:30.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-06-30" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:09.57">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-08-06" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:33.57">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-06-29" nation="" />
     <ATHLETE firstname="Carlo" nameprefix="" lastname="Travaini" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:27.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-06-04" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Emerson" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:02.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:23.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:21.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2014-08-17" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:08.20">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2014-08-15" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:29.36">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:01:03.60">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:02:19.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:04:54.43">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:10:32.07">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1958-11-25" />
    </RECORD>
    <RECORD swimtime="00:21:18.53">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-04" nation="NED" />
     <ATHLETE firstname="Donald" nameprefix="" lastname="Uijtenbogaart" gender="M" nation="NED" CLUB="Het Y" birthdate="1947-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:34.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Stockholm" date="2005-08-18" nation="SWE" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="De Veene" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:01:16.69">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2017-05-07" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:02:53.28">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:00:37.72">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Den Haag" date="2017-06-24" nation="NED" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Weyhenke" gender="M" nation="NED" CLUB="Upstream Amsterdam" birthdate="1952-07-29" />
    </RECORD>
    <RECORD swimtime="00:01:29.66">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2008-01-20" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="Neptunus" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:03:13.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Amsterdam" date="2008-10-25" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="Neptunus" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:00:29.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:01:05.82">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:32.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:02:38.68">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
    <RECORD swimtime="00:05:46.62">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Fukuoka" date="2023-08-07" nation="JPN" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" CLUB="WVZ" birthdate="1958-09-26" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:27.10">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Fukuoka" date="2023-08-09" nation="JPN" />
     <ATHLETE firstname="Igor" nameprefix="" lastname="Kravkov" gender="M" nation="ISR" />
    </RECORD>
    <RECORD swimtime="00:01:01.89">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2023-06-30" nation="ITA" />
     <ATHLETE firstname="Massimo" nameprefix="" lastname="Tubino" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:02:19.31">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Riccione" date="2023-06-29" nation="ITA" />
     <ATHLETE firstname="Massimo" nameprefix="" lastname="Tubino" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:04:54.43">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:10:13.58">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Villeurbanne" date="2022-04-30" nation="FRA" />
     <ATHLETE firstname="Serge" nameprefix="" lastname="Guerin" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:19:46.98">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Dijon" date="2023-05-13" nation="FRA" />
     <ATHLETE firstname="Serge" nameprefix="" lastname="Guerin" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:31.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Fukuoka" date="2023-08-11" nation="JPN" />
     <ATHLETE firstname="Igor" nameprefix="" lastname="Kravkov" gender="M" nation="ISR" />
    </RECORD>
    <RECORD swimtime="00:01:08.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="St. Petersburg" date="2022-04-22" nation="RUS" />
     <ATHLETE firstname="Vladimir" nameprefix="" lastname="Gorkov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:31.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="St. Petersburg" date="2022-04-23" nation="RUS" />
     <ATHLETE firstname="Vladimir" nameprefix="" lastname="Gorkov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:33.92">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Gwangju" date="2019-08-18" nation="KOR" />
     <ATHLETE firstname="Pere" nameprefix="" lastname="Balcells Prat" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:18.13">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Barcelona" date="2019-06-02" nation="ESP" />
     <ATHLETE firstname="Pere" nameprefix="" lastname="Balcells Prat" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:54.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Fukuoka" date="2023-08-10" nation="JPN" />
     <ATHLETE firstname="Sigitas" nameprefix="" lastname="Katkevicius" gender="M" nation="LTU" />
    </RECORD>
    <RECORD swimtime="00:00:28.54">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Girona" date="2009-06-27" nation="ESP" />
     <ATHLETE firstname="Josep" nameprefix="" lastname="Claret" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:05.82">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:32.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:38.68">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:05:42.24">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Pierrelatte" date="2018-06-30" nation="FRA" />
     <ATHLETE firstname="Patrick" nameprefix="" lastname="Moreau" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="65" agemax="69" />
   <RECORDS>
    <RECORD swimtime="00:00:26.21">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-07-06" nation="" />
     <ATHLETE firstname="Doug" nameprefix="" lastname="Martin" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:59.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-09-08" nation="" />
     <ATHLETE firstname="Jack" nameprefix="" lastname="Groselle" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:09.39">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-06" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:37.70">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-04" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:09:48.95">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-03" nation="" />
     <ATHLETE firstname="Djan" nameprefix="" lastname="Garrido Madruga" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:18:43.53">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-10-15" nation="" />
     <ATHLETE firstname="Paul" nameprefix="" lastname="Blackbeard" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:00:30.95">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2012-07-07" nation="" />
     <ATHLETE firstname="Hugh" nameprefix="" lastname="Wilder" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:08.15">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-04-22" nation="" />
     <ATHLETE firstname="Vladimir" nameprefix="" lastname="Gorkov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:02:31.62">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-04-23" nation="" />
     <ATHLETE firstname="Vladimir" nameprefix="" lastname="Gorkov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:33.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-08-19" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:14.77">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-08-05" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:41.54">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-08-21" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:28.26">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-07" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Thompson" gender="M" nation="CAN" />
    </RECORD>
    <RECORD swimtime="00:01:05.82">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:32.00">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
    </RECORD>
    <RECORD swimtime="00:02:25.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-08-19" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:13.36">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-08-03" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:31.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Harry" nameprefix="" lastname="Dokter" gender="M" nation="NED" CLUB="Swol 1894" birthdate="1951-07-04" />
    </RECORD>
    <RECORD swimtime="00:01:10.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:02:34.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Perth" date="2008-04-20" nation="AUS" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:05:33.24">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Perth" date="2008-04-24" nation="AUS" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:11:46.02">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Perth" date="2008-04-18" nation="AUS" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:23:33.45">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Luxembourg" date="2008-10-17" nation="LUX" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:00:36.43">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:01:21.27">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:03:02.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Antwerpen" date="2023-02-05" nation="BEL" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:00:40.64">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2008-01-19" nation="NED" />
     <ATHLETE firstname="Wieger" nameprefix="" lastname="Mensonides" gender="M" nation="NED" CLUB="NZ&amp;PC" birthdate="1938-07-12" />
    </RECORD>
    <RECORD swimtime="00:01:32.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-05-04" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:03:25.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-05-05" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:00:34.50">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" CLUB="PSV" birthdate="1952-02-26" />
    </RECORD>
    <RECORD swimtime="00:01:38.79">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Den Haag" date="2013-03-31" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:03:36.41">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Eindhoven" date="2013-09-04" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:03:09.88">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Perth" date="2008-04-21" nation="AUS" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Van Uden-de Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:07:10.36">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Wetzlar" date="2013-04-20" nation="GER" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:28.30">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Plymouth" date="2018-06-08" nation="GBR" />
     <ATHLETE firstname="John" nameprefix="" lastname="Liron" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:05.45">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2016-04-03" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:02:25.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2016-05-26" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:05:11.68">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2016-04-03" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:10:50.20">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Crawley" date="2016-01-23" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:21:05.22">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2017-03-04" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:34.81">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Elche" date="2016-02-21" nation="GER" />
     <ATHLETE firstname="Jean" nameprefix="" lastname="Lestideau" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:01:16.14">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2013-09-06" nation="NED" />
     <ATHLETE firstname="Bernd" nameprefix="" lastname="Horstmann" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:49.85">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2013-09-05" nation="NED" />
     <ATHLETE firstname="Bernd" nameprefix="" lastname="Horstmann" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:36.86">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kazan" date="2015-08-13" nation="RUS" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="H�fer" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:25.29">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-15" nation="HUN" />
     <ATHLETE firstname="Josef" nameprefix="" lastname="Kocsi" gender="M" nation="AUT" />
    </RECORD>
    <RECORD swimtime="00:03:11.63">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Josef" nameprefix="" lastname="Kocsi" gender="M" nation="AUT" />
    </RECORD>
    <RECORD swimtime="00:00:31.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Baltimore" date="2014-08-17" nation="USA" />
     <ATHLETE firstname="Josep" nameprefix="" lastname="Claret" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:14.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Montreal" date="2014-08-06" nation="CAN" />
     <ATHLETE firstname="Josep" nameprefix="" lastname="Claret" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:57.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Solingen" date="2022-03-20" nation="GER" />
     <ATHLETE firstname="Roland" nameprefix="" lastname="Freygang" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:51.06">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Antibes" date="2023-06-24" nation="FRA" />
     <ATHLETE firstname="Patrick" nameprefix="" lastname="Moreau" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:06:08.83">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Antibes" date="2023-06-23" nation="FRA" />
     <ATHLETE firstname="Patrick" nameprefix="" lastname="Moreau" gender="M" nation="FRA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="70" agemax="74" />
   <RECORDS>
    <RECORD swimtime="00:00:27.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-01-20" nation="USA" />
     <ATHLETE firstname="Doug" nameprefix="" lastname="Martin" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:03.32">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-08-08" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Quiggin" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:23.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-07-31" nation="" />
     <ATHLETE firstname="Fred" nameprefix="" lastname="Schlicher" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:57.84">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-07-01" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:10:12.57">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-07-01" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:20:26.12">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-07-20" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Kirkland" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:33.51">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-01-20" nation="USA" />
     <ATHLETE firstname="Bruce" nameprefix="" lastname="Williams" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:13.49">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-08-06" nation="" />
     <ATHLETE firstname="Hugh" nameprefix="" lastname="Wilder" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:40.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2021-06-05" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Day" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:34.69">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-07-01" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:17.80">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-07-01" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:48.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-07-01" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:29.98">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-10-10" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Day" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:07.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-10-08" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Day" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:47.17">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-10-09" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Day" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:35.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-07-01" nation="" />
     <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:55.97">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-06-06" nation="" />
     <ATHLETE firstname="Lawrence" nameprefix="" lastname="Day" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:33.33">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Apeldoorn" date="2001-06-16" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:17.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Munchen" date="2000-07-29" nation="GER" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:57.29">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kampen" date="2014-09-27" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Z&amp;PC De Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:06:22.00">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-09-02" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="Z&amp;PC De Gouwe" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:13:30.84">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Wout" nameprefix="" lastname="Hemmes" gender="M" nation="NED" CLUB="De Plons" birthdate="1948-06-16" />
    </RECORD>
    <RECORD swimtime="00:25:43.17">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-04" nation="NED" />
     <ATHLETE firstname="Wout" nameprefix="" lastname="Hemmes" gender="M" nation="NED" CLUB="De Plons" birthdate="1948-06-16" />
    </RECORD>
    <RECORD swimtime="00:00:38.57">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:01:25.84">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kazan" date="2015-08-15" nation="RUS" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:03:10.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kazan" date="2015-08-11" nation="RUS" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:00:42.76">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Eindhoven" date="2013-05-04" nation="NED" />
     <ATHLETE firstname="Wieger" nameprefix="" lastname="Mensonides" gender="M" nation="NED" CLUB="NZ&amp;PC" birthdate="1938-07-12" />
    </RECORD>
    <RECORD swimtime="00:01:36.52">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kranj" date="2018-09-07" nation="SLO" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:03:31.87">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kranj" date="2018-09-04" nation="SLO" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:00:40.03">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Kampen" date="2001-04-21" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:41.93">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Nijmegen" date="2001-05-26" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:04:50.67">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Copenhagen" date="2021-08-19" nation="DEN" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
    <RECORD swimtime="00:03:25.30">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Kazan" date="2015-08-13" nation="RUS" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:07:34.02">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Dordrecht" date="2019-02-17" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:30.11">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:01:09.37">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Dresden" date="2023-06-02" nation="GER" />
     <ATHLETE firstname="Dieter" nameprefix="" lastname="Seifert" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:35.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="London" date="2022-09-10" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:05:28.45">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Crawley" date="2023-01-21" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:11:24.63">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Crawley" date="2022-03-26" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:21:29.62">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Crawley" date="2022-03-26" nation="GBR" />
     <ATHLETE firstname="Christopher" nameprefix="" lastname="Dunn" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:00:36.32">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kranj" date="2018-09-07" nation="SLO" />
     <ATHLETE firstname="Jozsef" nameprefix="" lastname="Csikany" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:01:20.06">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kranj" date="2018-09-07" nation="SLO" />
     <ATHLETE firstname="Jozsef" nameprefix="" lastname="Csikany" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:58.32">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kranj" date="2018-09-06" nation="SLO" />
     <ATHLETE firstname="Jozsef" nameprefix="" lastname="Csikany" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:00:38.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Roma" date="2022-09-02" nation="ITA" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Rugieri" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:29.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Hannover" date="2011-07-01" nation="GER" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Reichelt" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:23.32">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Antibes" date="2023-06-22" nation="FRA" />
     <ATHLETE firstname="Alain" nameprefix="" lastname="Legrux" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:00:33.17">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Gwangju" date="2019-08-14" nation="KOR" />
     <ATHLETE firstname="Josep" nameprefix="" lastname="Claret" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:21.90">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Berlin" date="2022-03-13" nation="GER" />
     <ATHLETE firstname="Horst" nameprefix="" lastname="Lehmann" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:18.09">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Gwangju" date="2019-08-17" nation="KOR" />
     <ATHLETE firstname="Rudolf" nameprefix="" lastname="Smerda" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:03:03.47">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Roma" date="2022-08-31" nation="ITA" />
     <ATHLETE firstname="Josef" nameprefix="" lastname="Kocsi" gender="M" nation="AUT" />
    </RECORD>
    <RECORD swimtime="00:06:50.66">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Roma" date="2022-08-30" nation="ITA" />
     <ATHLETE firstname="Kurt" nameprefix="" lastname="Frei" gender="M" nation="SUI" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="75" agemax="79" />
   <RECORDS>
    <RECORD swimtime="00:00:29.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-08-25" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Quiggin" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:06.40">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-03-03" nation="" />
     <ATHLETE firstname="Akira" nameprefix="" lastname="Fujimaki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:25.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-06-06" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:17.77">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2009-03-07" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:11:01.70">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-11" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Kirkland" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:21:02.80">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-11" nation="" />
     <ATHLETE firstname="Dan" nameprefix="" lastname="Kirkland" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:34.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-08-02" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:17.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-07-31" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:50.25">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-07-30" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:38.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2022-09-02" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Rugieri" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:01:27.74">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-08-18" nation="" />
     <ATHLETE firstname="Mike" nameprefix="" lastname="Freshley" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:13.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2016-08-21" nation="" />
     <ATHLETE firstname="Mike" nameprefix="" lastname="Freshley" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:31.75">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-08-21" nation="" />
     <ATHLETE firstname="Joel" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:16.87">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-07-23" nation="" />
     <ATHLETE firstname="Fred" nameprefix="" lastname="Schlicher" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:08.54">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-07-22" nation="" />
     <ATHLETE firstname="Fred" nameprefix="" lastname="Schlicher" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:53.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-07-23" nation="" />
     <ATHLETE firstname="Joel" nameprefix="" lastname="Wilson" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:06:34.91">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-08-05" nation="" />
     <ATHLETE firstname="Mike" nameprefix="" lastname="Freshley" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:34.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Drachten" date="2004-01-24" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:21.86">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Drachten" date="2004-01-25" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:03:31.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="G�za" nameprefix="" lastname="Kaltenecker" gender="M" nation="NED" CLUB="AZC" birthdate="1942-10-20" />
    </RECORD>
    <RECORD swimtime="00:07:41.33">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <ATHLETE firstname="G�za" nameprefix="" lastname="Kaltenecker" gender="M" nation="NED" CLUB="AZC" birthdate="1942-10-20" />
    </RECORD>
    <RECORD swimtime="00:15:45.21">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-05" nation="NED" />
     <ATHLETE firstname="G�za" nameprefix="" lastname="Kaltenecker" gender="M" nation="NED" CLUB="AZC" birthdate="1942-10-20" />
    </RECORD>
    <RECORD swimtime="00:29:37.39">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-05" nation="NED" />
     <ATHLETE firstname="G�za" nameprefix="" lastname="Kaltenecker" gender="M" nation="NED" CLUB="AZC" birthdate="1942-10-20" />
    </RECORD>
    <RECORD swimtime="00:00:43.34">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Drachten" date="2004-01-24" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:40.21">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:03:39.38">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <ATHLETE firstname="Frans" nameprefix="van" lastname="Enst" gender="M" nation="NED" CLUB="WS Twente" birthdate="1940-02-01" />
    </RECORD>
    <RECORD swimtime="00:00:45.45">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kampen" date="2004-04-24" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:47.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Riccione" date="2004-06-07" nation="ITA" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:03:58.49">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kampen" date="2004-04-24" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:00:41.36">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Drachten" date="2004-01-25" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:49.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Riccione" date="2004-06-06" nation="ITA" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:03:44.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Riccione" date="2004-06-03" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:09:39.61">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" CLUB="PSV" birthdate="1943-12-25" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:31.28">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Kamen" date="2019-06-23" nation="GER" />
     <ATHLETE firstname="Helmut" nameprefix="" lastname="Richter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:13.12">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Las Palmas" date="2011-07-02" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:02:48.61">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gera" date="2016-04-16" nation="GER" />
     <ATHLETE firstname="Werner" nameprefix="" lastname="Schnabel" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:06:05.49">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Braunschweig" date="2016-02-28" nation="GER" />
     <ATHLETE firstname="Werner" nameprefix="" lastname="Schnabel" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:12:52.38">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Brescia" date="2011-03-06" nation="ITA" />
     <ATHLETE firstname="Giulio" nameprefix="" lastname="Divano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:24:40.69">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Genova" date="2011-05-15" nation="ITA" />
     <ATHLETE firstname="Giulio" nameprefix="" lastname="Divano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:39.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Szenes" date="2023-01-28" nation="HUN" />
     <ATHLETE firstname="Jozsef" nameprefix="" lastname="Csikany" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:01:26.31">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kecskemet" date="2023-04-15" nation="HUN" />
     <ATHLETE firstname="Jozsef" nameprefix="" lastname="Csikany" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:03:11.43">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Szentes" date="2023-01-28" nation="HUN" />
     <ATHLETE firstname="Jozsef" nameprefix="" lastname="Csikany" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:00:42.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-20" nation="HUN" />
     <ATHLETE firstname="Mikhail" nameprefix="" lastname="Farafonov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:34.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-15" nation="HUN" />
     <ATHLETE firstname="Bela" nameprefix="" lastname="Fabian" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:03:38.92">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-19" nation="HUN" />
     <ATHLETE firstname="Bela" nameprefix="" lastname="Fabian" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:00:36.73">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Pardubice" date="2023-04-22" nation="CZE" />
     <ATHLETE firstname="Rudolf" nameprefix="" lastname="Smerda" gender="M" nation="CZE" />
    </RECORD>
    <RECORD swimtime="00:01:29.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Brescia" date="2011-03-06" nation="ITA" />
     <ATHLETE firstname="Giulio" nameprefix="" lastname="Divano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:03:31.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2011-06-22" nation="ITA" />
     <ATHLETE firstname="Giulio" nameprefix="" lastname="Divano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:03:21.37">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Fukuoka" date="2023-08-08" nation="JPN" />
     <ATHLETE firstname="Gershon" nameprefix="" lastname="Shefa" gender="M" nation="ISR" />
    </RECORD>
    <RECORD swimtime="00:07:12.63">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Roma" date="2011-06-23" nation="ITA" />
     <ATHLETE firstname="Giulio" nameprefix="" lastname="Divano" gender="M" nation="ITA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="80" agemax="84" />
   <RECORDS>
    <RECORD swimtime="00:00:31.23">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-03-12" nation="" />
     <ATHLETE firstname="Akira" nameprefix="" lastname="Fujimaki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:08.76">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-03-11" nation="" />
     <ATHLETE firstname="Akira" nameprefix="" lastname="Fujimaki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:40.22">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-08-24" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:45.21">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2015-08-23" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:11:49.29">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-08-22" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:22:16.90">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2014-05-31" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:36.83">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-08-04" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:22.06">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-08-04" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:03:04.59">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2023-08-06" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:41.68">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2006-09-18" nation="" />
     <ATHLETE firstname="Toshio" nameprefix="" lastname="Tajima" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:34.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-08-01" nation="" />
     <ATHLETE firstname="Masaru" nameprefix="" lastname="Shinkai" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:27.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2021-08-01" nation="JPN" />
     <ATHLETE firstname="Masaru" nameprefix="" lastname="Shinkai" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:34.39">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-04" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:29.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2011-03-06" nation="" />
     <ATHLETE firstname="Divano" nameprefix="" lastname="Giulio" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:03:31.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Roma" date="2011-06-22" nation="ITA" />
     <ATHLETE firstname="Giulio" nameprefix="" lastname="Divano" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:03:15.52">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-06-17" nation="" />
     <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:07:12.03">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-10-24" nation="" />
     <ATHLETE firstname="Masaru" nameprefix="" lastname="Shinkai" gender="M" nation="JPN" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:42.81">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:01:37.69">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:03:51.93">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:08:38.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Alkmaar" date="2023-04-02" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:18:28.24">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-03" nation="NED" />
     <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" CLUB="PSV" birthdate="1933-04-17" />
    </RECORD>
    <RECORD swimtime="00:34:59.83">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-04" nation="NED" />
     <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" CLUB="PSV" birthdate="1938-07-24" />
    </RECORD>
    <RECORD swimtime="00:00:56.84">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2010-05-08" nation="NED" />
     <ATHLETE firstname="Ru" nameprefix="" lastname="Holtes" gender="M" nation="NED" CLUB="De Dolfijn" birthdate="1925-06-05" />
    </RECORD>
    <RECORD swimtime="00:01:58.55">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Cadiz" date="2009-09-19" nation="ESP" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:04:28.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Eindhoven" date="2010-05-07" nation="NED" />
     <ATHLETE firstname="Ru" nameprefix="" lastname="Holtes" gender="M" nation="NED" CLUB="De Dolfijn" birthdate="1925-06-05" />
    </RECORD>
    <RECORD swimtime="00:01:05.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Cadiz" date="2009-09-17" nation="ESP" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:12.92">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Apeldoorn" date="2009-06-13" nation="NED" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:01.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Cadiz" date="2009-09-15" nation="ESP" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="00:02:12.47">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Cadiz" date="2009-09-16" nation="ESP" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:04:29.94">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Cadiz" date="2009-09-15" nation="ESP" />
     <ATHLETE firstname="Max" nameprefix="van" lastname="Gelder" gender="M" nation="NED" CLUB="HZ&amp;PC Heerenveen" birthdate="1924-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:32.51">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Badajoz" date="2017-07-01" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:25.38">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Braunschweig" date="2021-09-10" nation="GER" />
     <ATHLETE firstname="Werner" nameprefix="" lastname="Schnabel" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:03.50">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Badajoz" date="2017-07-01" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:06:56.89">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Barcelona" date="2023-06-03" nation="ESP" />
     <ATHLETE firstname="Frederik-Henrik" nameprefix="" lastname="De Bruijn" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:14:18.23">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Barcelona" date="2023-04-29" nation="ESP" />
     <ATHLETE firstname="Frederik-Henrik" nameprefix="" lastname="De Bruijn" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:27:47.91">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Barcelona" date="2023-04-23" nation="ESP" />
     <ATHLETE firstname="Frederik-Henrik" nameprefix="" lastname="De Bruijn" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:00:45.58">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Badajoz" date="2017-07-01" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:42.86">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kranj" date="2018-09-04" nation="SLO" />
     <ATHLETE firstname="Fritz" nameprefix="" lastname="Ilgen" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:51.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kranj" date="2018-09-06" nation="SLO" />
     <ATHLETE firstname="Fritz" nameprefix="" lastname="Ilgen" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:46.08">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="St. Petersburg" date="2022-04-24" nation="RUS" />
     <ATHLETE firstname="Mikhail" nameprefix="" lastname="Farafonov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:01:46.19">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="San Francisco" date="2021-06-19" nation="USA" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Reichelt" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:03:58.36">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Mulhouse" date="2021-07-10" nation="FRA" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Reichelt" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:43.62">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Badajoz" date="2017-07-01" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:56.16">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-08" nation="JPN" />
     <ATHLETE firstname="David" nameprefix="" lastname="Cumming" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:04:14.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Fukuoka" date="2023-08-10" nation="JPN" />
     <ATHLETE firstname="David" nameprefix="" lastname="Cumming" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:57.74">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="G�teborg" date="2010-08-03" nation="SWE" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:08:34.82">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="K�ln" date="2010-04-23" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="85" agemax="89" />
   <RECORDS>
    <RECORD swimtime="00:00:33.74">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-08" nation="" />
     <ATHLETE firstname="Tohru" nameprefix="" lastname="Furukawa" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:22.25">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-08-06" nation="" />
     <ATHLETE firstname="Tohru" nameprefix="" lastname="Furukawa" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:03.50">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-07-01" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:06:38.87">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2016-06-26" nation="" />
     <ATHLETE firstname="Graham" nameprefix="" lastname="Johnston" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:13:56.29">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-07-19" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:26:18.37">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2019-07-19" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:39.89">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2008-07-18" nation="" />
     <ATHLETE firstname="Keijiro" nameprefix="" lastname="Nakamura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:31.65">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2008-03-02" nation="" />
     <ATHLETE firstname="Keijiro" nameprefix="" lastname="Nakamura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:03:28.59">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2008-07-19" nation="" />
     <ATHLETE firstname="Keijiro" nameprefix="" lastname="Nakamura" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:45.42">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-08-11" nation="" />
     <ATHLETE firstname="Tony" nameprefix="" lastname="Goodwin" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:01:40.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-08-06" nation="" />
     <ATHLETE firstname="Tony" nameprefix="" lastname="Goodwin" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:03:45.32">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2023-08-10" nation="" />
     <ATHLETE firstname="Tony" nameprefix="" lastname="Goodwin" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:00:43.62">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2017-07-01" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:50.27">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2021-04-11" nation="" />
     <ATHLETE firstname="John" nameprefix="" lastname="Cocks" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:04:14.19">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2023-08-10" nation="" />
     <ATHLETE firstname="David" nameprefix="" lastname="Cumming" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:39.66">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-03-21" nation="" />
     <ATHLETE firstname="John" nameprefix="" lastname="Cocks" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:07:56.23">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-03-20" nation="" />
     <ATHLETE firstname="John" nameprefix="" lastname="Cocks" gender="M" nation="AUS" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:01:13.39">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="00:03:05.39">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:04.29">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Alkmaar" date="2015-04-19" nation="NED" />
     <ATHLETE firstname="Ru" nameprefix="" lastname="Holtes" gender="M" nation="NED" CLUB="De Dolfijn" birthdate="1925-06-05" />
    </RECORD>
    <RECORD swimtime="00:03:14.41">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="00:01:52.51">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="00:04:10.43">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <ATHLETE firstname="Klaas" nameprefix="" lastname="Prins" gender="M" nation="NED" CLUB="Steenwijk 1934" birthdate="1928-08-10" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:00:38.64">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Murcia" date="2023-06-25" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:33.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Murcia" date="2023-06-24" nation="ESP" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:03:39.15">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Gera" date="2016-04-16" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:08:05.10">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Bari" date="2017-04-30" nation="ITA" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:17:29.90">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Wetzlar" date="2017-04-28" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:34:48.90">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="Scanzano Ionicoi" date="2017-05-27" nation="ITA" />
     <ATHLETE firstname="Domenic Antonio" nameprefix="" lastname="Casolino" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:00:51.01">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Braunschweig" date="2019-03-16" nation="GER" />
     <ATHLETE firstname="Karl-Heinz" nameprefix="" lastname="Klaustermeyer" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:01:58.06">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Fukuoka" date="2023-08-10" nation="JPN" />
     <ATHLETE firstname="Fritz" nameprefix="" lastname="Ilgen" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:17.01">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Aqua City" date="2023-09-23" nation="RUS" />
     <ATHLETE firstname="Valentin" nameprefix="" lastname="Meshcheryakov" gender="M" nation="RUS" />
    </RECORD>
    <RECORD swimtime="00:00:55.52">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Gera" date="2016-04-16" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:05.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Regensburg" date="2015-06-05" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:41.26">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Wetzlar" date="2017-04-30" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:54.13">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="Berlin" date="2022-03-12" nation="GER" />
     <ATHLETE firstname="Curt" nameprefix="" lastname="Zeiss" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:38.92">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="Regensburg" date="2015-06-06" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:06:05.42">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="Trieste" date="2005-07-08" nation="ITA" />
     <ATHLETE firstname="Aldo" nameprefix="" lastname="Caputi" gender="M" nation="ITA" />
    </RECORD>
    <RECORD swimtime="00:04:27.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="Regensburg" date="2015-06-05" nation="GER" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="90" agemax="94" />
   <RECORDS>
    <RECORD swimtime="00:00:38.64">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-06-24" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:01:33.00">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2023-06-24" nation="" />
     <ATHLETE firstname="Roberto" nameprefix="" lastname="Alberiche" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:03:33.64">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-12-12" nation="" />
     <ATHLETE firstname="Katsura" nameprefix="" lastname="Suzuki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:07:38.88">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-10-02" nation="" />
     <ATHLETE firstname="Katsura" nameprefix="" lastname="Suzuki" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:15:20.31">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-23" nation="" />
     <ATHLETE firstname="Katsuko" nameprefix="" lastname="Matsumoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:30:31.69">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2021-10-24" nation="" />
     <ATHLETE firstname="Katsuko" nameprefix="" lastname="Matsumoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:46.82">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2006-07-17" nation="" />
     <ATHLETE firstname="Goro" nameprefix="" lastname="Kobayashi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:01:45.46">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2006-08-09" nation="" />
     <ATHLETE firstname="Goro" nameprefix="" lastname="Kobayashi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:04:05.77">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2007-07-16" nation="" />
     <ATHLETE firstname="Goro" nameprefix="" lastname="Kobayashi" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:00:50.71">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2015-09-13" nation="" />
     <ATHLETE firstname="Toshio" nameprefix="" lastname="Tajima" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:05.18">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2015-06-05" nation="" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:04:41.26">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2017-04-30" nation="" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:00:54.13">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2022-03-12" nation="" />
     <ATHLETE firstname="Curt" nameprefix="" lastname="Zeiss" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:02:23.56">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2015-06-06" nation="" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Maine" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:19.18">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2015-06-06" nation="" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Maine" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:27.72">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-06-05" nation="" />
     <ATHLETE firstname="Karl" nameprefix="" lastname="Hauter" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="00:09:56.43">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-06-06" nation="" />
     <ATHLETE firstname="Thomas" nameprefix="" lastname="Maine" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:01:04.37">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Warszawa" date="2017-06-16" nation="POL" />
     <ATHLETE firstname="Kazimierz" nameprefix="" lastname="Mrowczynski" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:02:35.95">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-15" nation="HUN" />
     <ATHLETE firstname="Kazimierz" nameprefix="" lastname="Mrowczynski" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:05:36.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="Warszawa" date="2017-06-17" nation="POL" />
     <ATHLETE firstname="Kazimierz" nameprefix="" lastname="Mrowczynski" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:11:46.98">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="Mataro" date="2022-04-24" nation="ESP" />
     <ATHLETE firstname="Juan" nameprefix="" lastname="Dominguez" gender="M" nation="ESP" />
    </RECORD>
    <RECORD swimtime="00:22:07.69">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="Swansea" date="2023-03-05" nation="GBR" />
     <ATHLETE firstname="Edward" nameprefix="" lastname="Hoy" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="00:01:02.35">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kazan" date="2015-08-16" nation="RUS" />
     <ATHLETE firstname="Bela Banki" nameprefix="" lastname="Horvath" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:02:32.01">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kazan" date="2015-08-15" nation="RUS" />
     <ATHLETE firstname="Bela Banki" nameprefix="" lastname="Horvath" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:05:24.20">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="Kazan" date="2015-08-11" nation="RUS" />
     <ATHLETE firstname="Bela Banki" nameprefix="" lastname="Horvath" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:01:17.55">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-20" nation="HUN" />
     <ATHLETE firstname="Kazimierz" nameprefix="" lastname="Mrowczynski" gender="M" nation="POL" />
    </RECORD>
    <RECORD swimtime="00:04:39.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Budapest" date="2017-08-15" nation="HUN" />
     <ATHLETE firstname="Bela Banki" nameprefix="" lastname="Horvath" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="00:07:29.12">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="Kazan" date="2015-08-15" nation="RUS" />
     <ATHLETE firstname="Bela Banki" nameprefix="" lastname="Horvath" gender="M" nation="HUN" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="95" agemax="99" />
   <RECORDS>
    <RECORD swimtime="00:00:45.71">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-06" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:47.59">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-26" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:04.60">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-26" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:43.18">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-25" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:42.57">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-25" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:33:39.77">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2017-08-25" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:00:55.90">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2019-04-14" nation="" />
     <ATHLETE firstname="Anton" nameprefix="" lastname="Biedermann" gender="M" nation="BRA" />
    </RECORD>
    <RECORD swimtime="00:02:11.19">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2017-08-06" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:34.73">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2018-07-30" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:10.05">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2013-05-18" nation="" />
     <ATHLETE firstname="George" nameprefix="" lastname="Corones" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:02:40.08">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-06-20" nation="" />
     <ATHLETE firstname="Himoru" nameprefix="" lastname="Yoshimoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:05:47.31">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="2010-06-20" nation="" />
     <ATHLETE firstname="Himoru" nameprefix="" lastname="Yoshimoto" gender="M" nation="JPN" />
    </RECORD>
    <RECORD swimtime="00:02:01.41">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2008-06-01" nation="" />
     <ATHLETE firstname="Walter" nameprefix="" lastname="Pfeiffer" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:04:09.52">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2008-06-01" nation="" />
     <ATHLETE firstname="Walter" nameprefix="" lastname="Pfeiffer" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:11:47.68">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="2018-08-23" nation="" />
     <ATHLETE firstname="Robert" nameprefix="" lastname="Doud" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:08:55.97">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2008-06-01" nation="" />
     <ATHLETE firstname="Walter" nameprefix="" lastname="Pfeiffer" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:17:29.20">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="2008-06-01" nation="" />
     <ATHLETE firstname="Walter" nameprefix="" lastname="Pfeiffer" gender="M" nation="USA" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" CLUB="" birthdate="1900-01-01" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="00:01:31.19">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="Crawley" date="2014-02-01" nation="GBR" />
     <ATHLETE firstname="John" nameprefix="" lastname="Harrison" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="00:03:23.10">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="Crawley" date="2014-02-01" nation="GBR" />
     <ATHLETE firstname="John" nameprefix="" lastname="Harrison" gender="M" nation="GBR" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="00:01:29.13">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sarcelles" date="2014-05-04" nation="FRA" />
     <ATHLETE firstname="Jean" nameprefix="" lastname="Leemput" gender="M" nation="FRA" />
    </RECORD>
    <RECORD swimtime="00:06:01.50">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="Sindelfingen" date="2008-07-04" nation="GER" />
     <ATHLETE firstname="Hans" nameprefix="" lastname="Hahn" gender="M" nation="GER" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="104" />
   <RECORDS>
    <RECORD swimtime="00:00:56.12">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2018-02-28" nation="" />
     <ATHLETE firstname="George" nameprefix="" lastname="Corones" gender="M" nation="AUS" />
    </RECORD>
    <RECORD swimtime="00:02:15.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-07" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:18.86">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-03" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:10:55.25">
     <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-03" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:22:15.67">
     <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-03" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:42:27.06">
     <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
     <MEETINFO city="" date="2022-08-03" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:01:09.17">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-08-06" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:02:29.17">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2000-08-04" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="00:05:12.53">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
     <MEETINFO city="" date="2022-08-05" nation="" />
     <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="99" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:47.94">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <RELAY name="De Dolfijn" nation="NED">
      <CLUB name="De Dolfijn" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Tamara" nameprefix="" lastname="Grove" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Alinda" nameprefix="" lastname="Dingshoff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Romy" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Tessa" nameprefix="" lastname="Vermeulen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:01.92">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="STARTLIMIET" nation="">
      <CLUB name="STARTLIMIET" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:56.94">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-23" nation="NED" />
     <RELAY name="Aquarijn" nation="NED">
      <CLUB name="Aquarijn" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Linda" nameprefix="" lastname="Kamperman" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Richelle" nameprefix="" lastname="Koot" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Malissa" nameprefix="van der" lastname="Horst" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:28.06">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Terneuzen" date="2018-01-21" nation="NED" />
     <RELAY name="Hieronymus" nation="NED">
      <CLUB name="Hieronymus" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Eva" nameprefix="van" lastname="Ginneken" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Selene" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marlijn" nameprefix="" lastname="Hendriksen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nadja" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:57.06">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <RELAY name="Bubble" nation="NED">
      <CLUB name="Bubble" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Laura" nameprefix="" lastname="Setz" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Esmee" nameprefix="" lastname="Kloezen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marijke" nameprefix="" lastname="Drent" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Sanne" nameprefix="" lastname="Kloezen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:49.61">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Vlissingen" date="2005-03-06" nation="NED" />
     <RELAY name="SBC2000" nation="NED">
      <CLUB name="SBC2000" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Goossens" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Patricia" nameprefix="" lastname="Brooijmans" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Maartje" nameprefix="van" lastname="Keulen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Sandra" nameprefix="" lastname="Temmerman" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:56.42">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Britta" nameprefix="" lastname="Koehorst" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Anne Louise" nameprefix="" lastname="Palmans" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:00.03">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="Nuenen" nation="NED">
      <CLUB name="Nuenen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Richenne" nameprefix="" lastname="Zeebregts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Nikita" nameprefix="van den" lastname="Ouden" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Susan" nameprefix="" lastname="Teijken" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Anneloes" nameprefix="" lastname="Peulen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:24.86">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2015-01-24" nation="NED" />
     <RELAY name="De Dinkel" nation="NED">
      <CLUB name="De Dinkel" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Silke" nameprefix="" lastname="Oude Weernink" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Karin" nameprefix="" lastname="Hidding" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anique" nameprefix="" lastname="Willeme" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marlies" nameprefix="" lastname="Reinders" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:00.04">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <RELAY name="De Warande" nation="NED">
      <CLUB name="De Warande" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Amy" nameprefix="van" lastname="Lier" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Pauline" nameprefix="" lastname="Tieleman" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="D�sir�e" nameprefix="" lastname="Emmen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Melissa" nameprefix="van der" lastname="Geld" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:48.38">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="St. Petersburg" date="2015-11-29" nation="RUS" />
     <RELAY name="Neva Stars" nation="RUS">
      <CLUB name="Neva Stars" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:01.43">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Castellon" date="2023-02-19" nation="ESP" />
     <RELAY name="CN Monteverde" nation="ESP">
      <CLUB name="CN Monteverde" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:57.06">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Palma de Mallorca" date="2024-01-13" nation="ESP" />
     <RELAY name="Swim Camp Getxo" nation="ESP">
      <CLUB name="Swim Camp Getxo" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:24.86">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2015-01-24" nation="NED" />
     <RELAY name="De Dinkel" nation="NED">
      <CLUB name="De Dinkel" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Silke" nameprefix="" lastname="Oude Weernink" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Karin" nameprefix="" lastname="Hidding" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anique" nameprefix="" lastname="Willeme" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marlies" nameprefix="" lastname="Reinders" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:53.34">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2017-10-28" nation="GBR" />
     <RELAY name="Silver City" nation="GBR">
      <CLUB name="Silver City" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:45.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-05-21" nation="" />
     <RELAY name="Queendom" nation="JPN">
      <CLUB name="Queendom" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:54.05">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-05-21" nation="" />
     <RELAY name="Queendom" nation="JPN">
      <CLUB name="Queendom" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:55.76">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-11-17" nation="" />
     <RELAY name="SEN-SWIM" nation="JPN">
      <CLUB name="SEN-SWIM" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rie" nameprefix="" lastname="Nakagami" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kanako" nameprefix="" lastname="Tayama" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Maya" nameprefix="" lastname="Hatanaka" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Mika" nameprefix="" lastname="Kashiwazaki" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:14.24">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-09-23" nation="" />
     <RELAY name="RENAISSANCE" nation="JPN">
      <CLUB name="RENAISSANCE" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ayumi" nameprefix="" lastname="Watanabe" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Yoko" nameprefix="" lastname="Yamaguchi" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Mio" nameprefix="" lastname="Hirano" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Maki" nameprefix="" lastname="Mita" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:53.34">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-10-28" nation="" />
     <RELAY name="SILVER CITY" nation="GBR">
      <CLUB name="SILVER CITY" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rachael" nameprefix="" lastname="Keir" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Louise" nameprefix="" lastname="Kennedy" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Kelly" nameprefix="" lastname="Mcintosh" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Laura" nameprefix="" lastname="Robertson" gender="F" nation="GBR" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:50.88">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zuidbroek" date="2003-11-15" nation="NED" />
     <RELAY name="AZ&amp;PC" nation="NED">
      <CLUB name="AZ&amp;PC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Tamara" nameprefix="van" lastname="Gorkom" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:05.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lauren" nameprefix="van" lastname="IJll" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Manon" nameprefix="van" lastname="Strien" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:06.40">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lauren" nameprefix="van" lastname="IJll" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Manon" nameprefix="van" lastname="Strien" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:38.67">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Manon" nameprefix="van" lastname="Strien" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lauren" nameprefix="van" lastname="IJll" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:20.10">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-24" nation="NED" />
     <RELAY name="Het Y" nation="NED">
      <CLUB name="Het Y" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Bravo" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Cynthia" nameprefix="" lastname="Noordermeer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ana-Lara" nameprefix="da" lastname="Silva" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Evelien" nameprefix="" lastname="Sohl" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:44.88">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="St. Petersburg" date="2014-11-30" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novgorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novgorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:56.67">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Risenga" date="2008-03-06" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novgorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novgorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:56.12">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Antwerpen" date="2021-12-17" nation="BEL" />
     <RELAY name="Brabo Antwerpen" nation="BEL">
      <CLUB name="Brabo Antwerpen" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:24.80">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2017-10-28" nation="GBR" />
     <RELAY name="Teddington Masters" nation="GBR">
      <CLUB name="Teddington Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:50.47">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2018-10-27" nation="GBR" />
     <RELAY name="Teddington Masters" nation="GBR">
      <CLUB name="Teddington Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:44.88">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2014-11-30" nation="" />
     <RELAY name="TSUNAMI" nation="RUS">
      <CLUB name="TSUNAMI" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Irina" nameprefix="" lastname="Shlemova" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Liubov" nameprefix="" lastname="Yudina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ekatarina" nameprefix="" lastname="Yudina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Svetlana" nameprefix="" lastname="Kniaginina" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:54.21">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-04-17" nation="" />
     <RELAY name="Team Go Mai Way" nation="JPN">
      <CLUB name="Team Go Mai Way" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:56.12">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-12-17" nation="" />
     <RELAY name="Brabo" nation="BEL">
      <CLUB name="Brabo" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:24.80">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-10-28" nation="" />
     <RELAY name="TEDDINSTON MASTERS" nation="GBR">
      <CLUB name="TEDDINSTON MASTERS" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Hannah" nameprefix="" lastname="Loughlin" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Georgina" nameprefix="" lastname="Heyn" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rebecca" nameprefix="" lastname="Newson" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Zoe" nameprefix="" lastname="Liokalos" gender="F" nation="GBR" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:42.32">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-12-03" nation="" />
     <RELAY name="TNT/Okuda" nation="BRA">
      <CLUB name="TNT/Okuda" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:53.16">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2004-02-21" nation="NED" />
     <RELAY name="AZ&amp;PC " nation="NED">
      <CLUB name="AZ&amp;PC " nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Petra" nameprefix="" lastname="Casteleijn-Frowijn" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:09.39">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Steenwijk" date="2019-09-14" nation="NED" />
     <RELAY name="Zpc Amersfoort" nation="NED">
      <CLUB name="Zpc Amersfoort" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:15.85">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-12-03" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lisa" nameprefix="" lastname="Dreesens" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:39.06">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2016-12-03" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lisa" nameprefix="" lastname="Dreesens" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:40.49">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2009-10-31" nation="NED" />
     <RELAY name="AZ&amp;PC" nation="NED">
      <CLUB name="AZ&amp;PC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Fran�oise" nameprefix="" lastname="Duran" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:47.58">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Saransk" date="2019-11-24" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novgorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novgorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:00.84">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Helsingborg" date="2016-05-08" nation="SWE" />
     <RELAY name="Helsingborgs Sims�llskap" nation="SWE">
      <CLUB name="Helsingborgs Sims�llskap" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:02.15">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-27" nation="GBR" />
     <RELAY name="Basingstoke" nation="GBR">
      <CLUB name="Basingstoke" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:35.01">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2018-10-27" nation="GBR" />
     <RELAY name="Teddington Masters" nation="GBR">
      <CLUB name="Teddington Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:54.33">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-28" nation="GBR" />
     <RELAY name="Basingstoke" nation="GBR">
      <CLUB name="Basingstoke" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:47.58">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-11-24" nation="" />
     <RELAY name="TSUNAMI" nation="RUS">
      <CLUB name="TSUNAMI" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Irina" nameprefix="" lastname="Shlemova" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Liubov" nameprefix="" lastname="Yudina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ekatarina" nameprefix="" lastname="Yudina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Olga" nameprefix="" lastname="Borisova" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:59.33">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-03-18" nation="" />
     <RELAY name="North Carolina Masters" nation="USA">
      <CLUB name="North Carolina Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:02.15">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-10-27" nation="" />
     <RELAY name="Basingstoke" nation="GBR">
      <CLUB name="Basingstoke" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:31.32">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-11-17" nation="" />
     <RELAY name="NORTH CAROLINA MASTERS" nation="USA">
      <CLUB name="NORTH CAROLINA MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kerry" nameprefix="" lastname="Lindauer" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Sarah" nameprefix="" lastname="Dunn" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Irish" nameprefix="" lastname="Holland" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:54.33">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-10-28" nation="" />
     <RELAY name="Basingstoke" nation="GBR">
      <CLUB name="Basingstoke" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:56.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:13.08">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jeanne" nameprefix="" lastname="Petit" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:18.18">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:50.03">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jeanne" nameprefix="" lastname="Petit" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:18.55">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:56.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:08.77">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Bergen" date="2019-03-08" nation="NOR" />
     <RELAY name="Masters Sorlandet" nation="NOR">
      <CLUB name="Masters Sorlandet" nation="NOR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:17.02">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Palma de Mallorca" date="2022-04-23" nation="ESP" />
     <RELAY name="T�r�kbalin" nation="HUN">
      <CLUB name="T�r�kbalin" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:50.03">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jeanne" nameprefix="" lastname="Petit" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:18.55">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:54.26">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2020-02-29" nation="" />
     <RELAY name="Club Tribe Alumn" nation="USA">
      <CLUB name="Club Tribe Alumn" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:06.51">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-12-04" nation="" />
     <RELAY name="Club Tribe" nation="USA">
      <CLUB name="Club Tribe" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:17.02">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-04-23" nation="" />
     <RELAY name="Torokbalin" nation="HUN">
      <CLUB name="Torokbalin" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:48.61">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-11-08" nation="" />
     <RELAY name="NORTH TEXAS MASTERS" nation="USA">
      <CLUB name="NORTH TEXAS MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Stephanie" nameprefix="" lastname="Stone" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Maureen" nameprefix="" lastname="Rea" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lisa" nameprefix="" lastname="Mize" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lynn" nameprefix="" lastname="Morrison" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:18.55">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:19.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Leiden" date="2023-09-17" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:26.24">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Krupiarz" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jeanne" nameprefix="" lastname="Petit" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:04.38">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2023-11-26" nation="NED" />
     <RELAY name="Psv" nation="NED">
      <CLUB name="Psv" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Katrin" nameprefix="" lastname="Pennings" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:48.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2023-11-26" nation="NED" />
     <RELAY name="Psv" nation="NED">
      <CLUB name="Psv" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:11:38.59">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <RELAY name="Swol 1894" nation="NED">
      <CLUB name="Swol 1894" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Bea" nameprefix="" lastname="Swijnenberg" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Mathilde" nameprefix="" lastname="Vink" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Annemarie" nameprefix="" lastname="Vuist-Blum" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:06.79">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2019-10-26" nation="GBR" />
     <RELAY name="Camp Hill Edwardians" nation="GBR">
      <CLUB name="Camp Hill Edwardians" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:20.46">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:51.67">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-27" nation="GBR" />
     <RELAY name="Gateshead &amp; Whickham" nation="GBR">
      <CLUB name="Gateshead &amp; Whickham" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:18.65">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:27.21">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2019-10-26" nation="GBR" />
     <RELAY name="Camphill Edwardians" nation="GBR">
      <CLUB name="Camphill Edwardians" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:02.15">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-11-11" nation="" />
     <RELAY name="NORTH TEXAS MASTERS" nation="USA">
      <CLUB name="NORTH TEXAS MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kristin" nameprefix="" lastname="Henderson" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lynn" nameprefix="" lastname="Morisson" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Christina" nameprefix="" lastname="Mckelvey" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Monica" nameprefix="" lastname="Bailey" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:18.67">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-10-07" nation="" />
     <RELAY name="Kana Kana" nation="JPN">
      <CLUB name="Kana Kana" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:30.74">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2016-03-06" nation="" />
     <RELAY name="UCLA" nation="USA">
      <CLUB name="UCLA" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jacki" nameprefix="" lastname="Hirsty" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Christie" nameprefix="" lastname="Ciraulo" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jenny" nameprefix="" lastname="Cook" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Veronica" nameprefix="" lastname="Hibben" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:07.72">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-03-11" nation="" />
     <RELAY name="Oregon Masters" nation="USA">
      <CLUB name="Oregon Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:09.82">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-10-13" nation="" />
     <RELAY name="Swim Melbourne" nation="AUS">
      <CLUB name="Swim Melbourne" nation="AUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:25.83">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Krupiarz" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:48.97">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:21.18">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:39.47">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Krupiarz" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:12:06.47">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:25.83">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Krupiarz" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:44.11">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Copenhagen" date="2023-11-04" nation="DEN" />
     <RELAY name="Swim Team Taastrup" nation="DEN">
      <CLUB name="Swim Team Taastrup" nation="DEN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:21.18">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:12.17">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <RELAY name="Spencer Swim Team" nation="GBR">
      <CLUB name="Spencer Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:12:06.47">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-25" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:14.25">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-01-21" nation="" />
     <RELAY name="Lone Star Masters" nation="USA">
      <CLUB name="Lone Star Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:32.54">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-01-22" nation="" />
     <RELAY name="Lone Star Masters" nation="USA">
      <CLUB name="Lone Star Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:03.06">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-01-22" nation="" />
     <RELAY name="Lone Star Masters" nation="USA">
      <CLUB name="Lone Star Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:54.73">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-01-21" nation="" />
     <RELAY name="Lone Star Masters" nation="USA">
      <CLUB name="Lone Star Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:11:54.09">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-10-14" nation="" />
     <RELAY name="Sarasota Sharks Masters" nation="USA">
      <CLUB name="Sarasota Sharks Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:04.54">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:54.89">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-12-03" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Annie" nameprefix="" lastname="Smits" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:25.40">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2016-12-03" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:03:05.64">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Helsingborg" date="2007-03-24" nation="SWE" />
     <RELAY name="SOIK HELLAS" nation="SWE">
      <CLUB name="SOIK HELLAS" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:52.52">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Helsingb�rg" date="2007-03-25" nation="SWE" />
     <RELAY name="Hellas Masters" nation="SWE">
      <CLUB name="Hellas Masters" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:51.31">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="London" date="2019-07-07" nation="GBR" />
     <RELAY name="Spencer Swim Team" nation="GBR">
      <CLUB name="Spencer Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:20.97">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="London" date="2019-07-07" nation="GBR" />
     <RELAY name="Spencer Swim Team" nation="GBR">
      <CLUB name="Spencer Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:17:13.93">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="London" date="2019-07-07" nation="GBR" />
     <RELAY name="Spencer Swim Team" nation="GBR">
      <CLUB name="Spencer Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:55.60">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2013-02-16" nation="" />
     <RELAY name="BIG S YOKOHAMA" nation="JPN">
      <CLUB name="BIG S YOKOHAMA" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Sonoe" nameprefix="" lastname="Watanabe" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Meiko" nameprefix="" lastname="Kamashita" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Masae" nameprefix="" lastname="Kurata" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:16.89">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-01-22" nation="" />
     <RELAY name="St Kansai" nation="JPN">
      <CLUB name="St Kansai" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:40.83">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-06-19" nation="" />
     <RELAY name="Miami Masters" nation="USA">
      <CLUB name="Miami Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:48.04">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-05-22" nation="" />
     <RELAY name="Miami Masters" nation="AUS">
      <CLUB name="Miami Masters" nation="AUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:16:13.28">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-10-21" nation="" />
     <RELAY name="SUNWAY YOKOHAMA" nation="JPN">
      <CLUB name="SUNWAY YOKOHAMA" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Sachie" nameprefix="" lastname="Mori" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Yuko" nameprefix="" lastname="Sakagami" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Sonoe" nameprefix="" lastname="Watanabe" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:04:45.07">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2013-06-02" nation="" />
     <RELAY name="SAPPORO MASTERS" nation="JPN">
      <CLUB name="SAPPORO MASTERS" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kinko" nameprefix="" lastname="Matsumoto" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Setsuko" nameprefix="" lastname="Narita" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Naka" nameprefix="" lastname="Fukuoka" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fumi" nameprefix="" lastname="Murata" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:40.08">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-03-06" nation="" />
     <RELAY name="SAPPORO MASTERS" nation="JPN">
      <CLUB name="SAPPORO MASTERS" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Sumiko" nameprefix="" lastname="Kuji" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Naka" nameprefix="" lastname="Fukuoka" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Haruko" nameprefix="" lastname="Sasaki" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fumi" nameprefix="" lastname="Murata" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="99" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:36.53">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-25" nation="NED" />
     <RELAY name="RZC" nation="NED">
      <CLUB name="RZC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Stefan" nameprefix="" lastname="Timmermans" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kevin" nameprefix="van" lastname="Susteren" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Raynor" nameprefix="" lastname="Wolf" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Pascal" nameprefix="" lastname="Timmermans" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:47.81">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Kuipers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Gavin" nameprefix="van der" lastname="Werf" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jorian" nameprefix="" lastname="Darwinkel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Remco" nameprefix="" lastname="Dijkstra" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:35.57">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="Albion WSS (SG)" nation="NED">
      <CLUB name="Albion WSS (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ayrton" nameprefix="" lastname="Mooldijk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Otto" nameprefix="" lastname="Pranger" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Pascal" nameprefix="" lastname="Nuijten" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:58.07">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Kuipers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Gavin" nameprefix="van der" lastname="Werf" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jorian" nameprefix="" lastname="Darwinkel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Remco" nameprefix="" lastname="Dijkstra" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:52.24">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <RELAY name="Albion WSS (SG)" nation="NED">
      <CLUB name="Albion WSS (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Thomas" nameprefix="" lastname="Verhoeven" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Pascal" nameprefix="" lastname="Nuijten" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:35.09">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="Rotterdam Swimming (SG)" nation="NED">
      <CLUB name="Rotterdam Swimming (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Derk Jan" nameprefix="" lastname="Speelman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Melvin" nameprefix="" lastname="Prins" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Martijn" nameprefix="" lastname="Dolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:48.57">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="De Kempvis" nation="NED">
      <CLUB name="De Kempvis" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Joris" nameprefix="" lastname="Bezemer" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Floyd" nameprefix="van" lastname="Duyvenbode" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Wegman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:31.31">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <RELAY name="Feijenoord Albion Zwemclub" nation="NED">
      <CLUB name="Feijenoord Albion Zwemclub" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:50.38">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <RELAY name="Feijenoord Albion Zwemclub" nation="NED">
      <CLUB name="Feijenoord Albion Zwemclub" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:10.47">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-24" nation="NED" />
     <RELAY name="ZPC DE HOF" nation="NED">
      <CLUB name="ZPC DE HOF" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Pieter" nameprefix="" lastname="Pickhardt" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jasper" nameprefix="de" lastname="Boer" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Emiel" nameprefix="" lastname="Huisken" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Huisken" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:31.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Kastrup" date="2009-11-07" nation="DEN" />
     <RELAY name="USG RACE CLUB" nation="DEN">
      <CLUB name="USG RACE CLUB" nation="DEN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:38.97">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Tallin" date="2021-09-25" nation="EST" />
     <RELAY name="Kalevi Ujumiskool" nation="EST">
      <CLUB name="Kalevi Ujumiskool" nation="EST" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:24.53">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2019-10-27" nation="GBR" />
     <RELAY name="East Leeds" nation="GBR">
      <CLUB name="East Leeds" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:41.62">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2023-10-27" nation="GBR" />
     <RELAY name="Dartmoor Dartes" nation="GBR">
      <CLUB name="Dartmoor Dartes" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:40.86">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Farum" date="2016-05-22" nation="DEN" />
     <RELAY name="Sarum Swommeklub" nation="DEN">
      <CLUB name="Sarum Swommeklub" nation="DEN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:30.73">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2009-12-12" nation="" />
     <RELAY name="OKUDINHAS" nation="BRA">
      <CLUB name="OKUDINHAS" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ricardo" nameprefix="" lastname="Wassall" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Daniel" nameprefix="" lastname="Belini" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Leandro" nameprefix="" lastname="Okuda" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Alexander" nameprefix="" lastname="Rehder" gender="M" nation="BRA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:38.97">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-09-25" nation="" />
     <RELAY name="Kalevi Ijumiskool" nation="EST">
      <CLUB name="Kalevi Ijumiskool" nation="EST" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:24.53">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-10-27" nation="" />
     <RELAY name="EAST LEEDS SWIM CLUB" nation="GBR">
      <CLUB name="EAST LEEDS SWIM CLUB" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Alistair" nameprefix="" lastname="Crawford" gender="M" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Jagger" gender="M" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Ayre" gender="M" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ryan" nameprefix="" lastname="Flanagan" gender="M" nation="GBR" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:41.62">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-10-27" nation="" />
     <RELAY name="Dartmoor Darts" nation="GBR">
      <CLUB name="Dartmoor Darts" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:18.39">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-05-16" nation="" />
     <RELAY name="JFE Keihin" nation="JPN">
      <CLUB name="JFE Keihin" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:35.70">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <RELAY name="Feijenoord Albion Zwemclub" nation="NED">
      <CLUB name="Feijenoord Albion Zwemclub" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Bart" nameprefix="" lastname="Drechsel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:46.28">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <RELAY name="Feijenoord Albion Zwemclub" nation="NED">
      <CLUB name="Feijenoord Albion Zwemclub" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Bart" nameprefix="" lastname="Drechsel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:35.42">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-23" nation="NED" />
     <RELAY name="d&apos;ELFT WAVE (SG)" nation="NED">
      <CLUB name="d&apos;ELFT WAVE (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Roderik" nameprefix="" lastname="Meijers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:59.37">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Papendrecht" date="2016-01-24" nation="NED" />
     <RELAY name="d&apos;ELFT WAVE (SG)" nation="NED">
      <CLUB name="d&apos;ELFT WAVE (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Roderik" nameprefix="" lastname="Meijers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:08.40">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <RELAY name="d&apos;ELFT WAVE (SG)" nation="NED">
      <CLUB name="d&apos;ELFT WAVE (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Roderik" nameprefix="" lastname="Meijers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:30.83">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Saransk" date="2019-11-24" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novgorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novgorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:43.56">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2009-10-24" nation="GBR" />
     <RELAY name="Swindon Dolphins" nation="GBR">
      <CLUB name="Swindon Dolphins" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:27.54">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Santurtzi" date="2014-05-10" nation="ESP" />
     <RELAY name="GETXO I.WP" nation="ESP">
      <CLUB name="GETXO I.WP" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:47.57">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <RELAY name="East Leeds" nation="GBR">
      <CLUB name="East Leeds" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:42.60">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Gussago" date="2017-01-29" nation="ITA" />
     <RELAY name="Brescia Acquare Mafeco" nation="ITA">
      <CLUB name="Brescia Acquare Mafeco" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:30.83">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-11-24" nation="" />
     <RELAY name="TSUNAMI" nation="RUS">
      <CLUB name="TSUNAMI" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Aleksey" nameprefix="" lastname="Getmanenko" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Alexandr" nameprefix="" lastname="Satanovskiy" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Sergey" nameprefix="" lastname="Mukhin" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Andrei" nameprefix="" lastname="Kurnosov" gender="M" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:38.46">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-03-18" nation="" />
     <RELAY name="JFE KEIHIN" nation="JPN">
      <CLUB name="JFE KEIHIN" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Takashi" nameprefix="" lastname="Takemoto" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Yuuki" nameprefix="" lastname="Kanaya" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ryoya" nameprefix="" lastname="Taguchi" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Shintaro" nameprefix="" lastname="Uchiyama" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:23.55">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2018-05-20" nation="" />
     <RELAY name="JFE KEIHIN" nation="JPN">
      <CLUB name="JFE KEIHIN" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ryoya" nameprefix="" lastname="Taguchi" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Takashi" nameprefix="" lastname="Takemoto" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Takao" nameprefix="" lastname="Ueki" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Shintaro" nameprefix="" lastname="Uchiyama" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:38.08">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-02-12" nation="" />
     <RELAY name="Diablo" nation="JPN">
      <CLUB name="Diablo" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:30.89">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-04-09" nation="" />
     <RELAY name="BLUE CORSAIRS" nation="JPN">
      <CLUB name="BLUE CORSAIRS" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ryoya" nameprefix="" lastname="Taguchi" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Takashi" nameprefix="" lastname="Takemoto" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Shintaro" nameprefix="" lastname="Uchiyama" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Takao" nameprefix="" lastname="Ueki" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:38.57">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Vincent" nameprefix="" lastname="Bakker" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Joan" nameprefix="" lastname="Kentrop" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:50.35">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <RELAY name="Albion d&apos;ELFT (SG)" nation="NED">
      <CLUB name="Albion d&apos;ELFT (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:39.90">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-21" nation="NED" />
     <RELAY name="Albion d&apos;ELFT (SG)" nation="NED">
      <CLUB name="Albion d&apos;ELFT (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:03.20">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <RELAY name="Albion d&apos;ELFT (SG)" nation="NED">
      <CLUB name="Albion d&apos;ELFT (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:15.42">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-20" nation="NED" />
     <RELAY name="Albion d&apos;ELFT (SG)" nation="NED">
      <CLUB name="Albion d&apos;ELFT (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:32.77">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Castellon" date="2023-02-18" nation="ESP" />
     <RELAY name="Swim camp Getxo CD" nation="ESP">
      <CLUB name="Swim camp Getxo CD" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:42.65">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Milano" date="2023-12-17" nation="ITA" />
     <RELAY name="Aquamore - Acqua 13" nation="ITA">
      <CLUB name="Aquamore - Acqua 13" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:27.42">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Mol" date="2019-03-23" nation="BEL" />
     <RELAY name="MOZKA" nation="BEL">
      <CLUB name="MOZKA" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:49.40">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Milano" date="2023-12-16" nation="ITA" />
     <RELAY name="Aquamore - Acqual 13" nation="ITA">
      <CLUB name="Aquamore - Acqual 13" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:52.68">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Glostrup" date="2016-03-12" nation="DEN" />
     <RELAY name="Sigma Swim" nation="DEN">
      <CLUB name="Sigma Swim" nation="DEN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:32.77">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-02-18" nation="" />
     <RELAY name="SC Getxo" nation="ESP">
      <CLUB name="SC Getxo" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:42.90">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-02-11" nation="" />
     <RELAY name="Diablo" nation="JPN">
      <CLUB name="Diablo" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:27.42">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-03-23" nation="" />
     <RELAY name="MOZKA" nation="BEL">
      <CLUB name="MOZKA" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Fr�d�ric" nameprefix="" lastname="Tonus" gender="M" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ruud" nameprefix="" lastname="Cuyvers" gender="M" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Michel" nameprefix="Van" lastname="Thielen" gender="M" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Stef" nameprefix="" lastname="Verachten" gender="M" nation="BEL" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:47.97">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-01-29" nation="" />
     <RELAY name="JSS Fukai" nation="JPN">
      <CLUB name="JSS Fukai" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:48.49">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-08-08" nation="" />
     <RELAY name="JSS Fukai" nation="JPN">
      <CLUB name="JSS Fukai" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:45.02">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <RELAY name="De Rog" nation="NED">
      <CLUB name="De Rog" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Spetter" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Arjan" nameprefix="" lastname="Verheij" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Glen" nameprefix="le" lastname="Clercq" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:56.95">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Joost" nameprefix="" lastname="Groeneveld" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Gijsbert" nameprefix="van der" lastname="Leden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:57.04">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-23" nation="NED" />
     <RELAY name="De Rog" nation="NED">
      <CLUB name="De Rog" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Spetter" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Kamphuis" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Glen" nameprefix="le" lastname="Clercq" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:25.59">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ivo" nameprefix="" lastname="Roozeboom" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jan-Willem" nameprefix="van den" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Markus" nameprefix="van" lastname="Rest" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:04.60">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Papendrecht" date="2016-01-22" nation="NED" />
     <RELAY name="De Rog" nation="NED">
      <CLUB name="De Rog" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Spetter" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Kamphuis" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Glen" nameprefix="le" lastname="Clercq" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:38.57">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Saransk" date="2021-11-14" nation="RUS" />
     <RELAY name="Mad Wave" nation="RUS">
      <CLUB name="Mad Wave" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:49.80">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2021-11-13" nation="RUS" />
     <RELAY name="Mad Wave" nation="RUS">
      <CLUB name="Mad Wave" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:39.17">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Gussago" date="2017-01-28" nation="ITA" />
     <RELAY name="Brescia Acquare Mafeco" nation="ITA">
      <CLUB name="Brescia Acquare Mafeco" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:13.39">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <RELAY name="Warrington Masters" nation="GBR">
      <CLUB name="Warrington Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:14.56">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <RELAY name="I.L. Varg" nation="NOR">
      <CLUB name="I.L. Varg" nation="NOR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jarl Inge" nameprefix="" lastname="Melberg" gender="M" nation="NOR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Oddvar" nameprefix="" lastname="Sandvin" gender="M" nation="NOR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="�ivind Martin" nameprefix="" lastname="Hasle" gender="M" nation="NOR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Erlend" nameprefix="" lastname="Alstad" gender="M" nation="NOR" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:37.35">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-05-28" nation="" />
     <RELAY name="Tattersalls Masters" nation="AUS">
      <CLUB name="Tattersalls Masters" nation="AUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:48.40">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-05-07" nation="" />
     <RELAY name="MTR" nation="JPN">
      <CLUB name="MTR" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:40.26">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2011-10-15" nation="" />
     <RELAY name="BLU FROG TEAM" nation="USA">
      <CLUB name="BLU FROG TEAM" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Charles" nameprefix="" lastname="Lydecker" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ross" nameprefix="" lastname="Bohlken" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Keith" nameprefix="" lastname="Switzer" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ambrose" nameprefix="" lastname="Gaines" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:59.68">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2012-12-02" nation="" />
     <RELAY name="LONGHORN AQUATICS" nation="USA">
      <CLUB name="LONGHORN AQUATICS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Anders" nameprefix="" lastname="Rasmussen" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jim" nameprefix="" lastname="Sauer" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="David" nameprefix="" lastname="Guthrie" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Mike" nameprefix="" lastname="Varozza" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:03.40">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2011-10-14" nation="" />
     <RELAY name="BLU FROG TEAM" nation="USA">
      <CLUB name="BLU FROG TEAM" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ambrose" nameprefix="" lastname="Gaines" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Charles" nameprefix="" lastname="Lydecker" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Tim" nameprefix="" lastname="Buckley" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Keith" nameprefix="" lastname="Switzer" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:52.33">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Joop" nameprefix="" lastname="Ariaens" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:07.37">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Evertjan" nameprefix="" lastname="Masurel" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:15.08">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Weert" date="2017-03-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Joop" nameprefix="" lastname="Ariaens" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:50.13">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Joop" nameprefix="" lastname="Ariaens" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:26.62">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-24" nation="NED" />
     <RELAY name="WWV Winterswijk" nation="NED">
      <CLUB name="WWV Winterswijk" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kees-Jan" nameprefix="van" lastname="Overbeeke" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Laurens" nameprefix="" lastname="Klein Breteler" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Theo" nameprefix="" lastname="Schouten" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ruud" nameprefix="" lastname="Ruiter" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:47.90">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Dunkerque" date="2017-03-23" nation="FRA" />
     <RELAY name="SF Coubevoie" nation="FRA">
      <CLUB name="SF Coubevoie" nation="FRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:00.94">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rennes" date="2015-03-28" nation="FRA" />
     <RELAY name="SFO Courbevoie" nation="FRA">
      <CLUB name="SFO Courbevoie" nation="FRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:10.69">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-27" nation="GBR" />
     <RELAY name="Warrender Baths" nation="GBR">
      <CLUB name="Warrender Baths" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:34.10">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Desenzano" date="2019-01-26" nation="ITA" />
     <RELAY name="Nuoto Master Brescia" nation="ITA">
      <CLUB name="Nuoto Master Brescia" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:18.30">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Saransk" date="2021-11-14" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novogorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novogorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:43.21">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2012-10-14" nation="" />
     <RELAY name="BLU FROG TEAM" nation="USA">
      <CLUB name="BLU FROG TEAM" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ambrose" nameprefix="" lastname="Gaines" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marc" nameprefix="" lastname="Middleton" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Keith" nameprefix="" lastname="Switzer" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Scot" nameprefix="" lastname="Weiss" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:54.15">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-11-10" nation="" />
     <RELAY name="RICE AQUATIC MASTERS" nation="USA">
      <CLUB name="RICE AQUATIC MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jay" nameprefix="" lastname="Yarid" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="David" nameprefix="" lastname="Guthrie" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="John" nameprefix="" lastname="Fields" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Bruce" nameprefix="" lastname="Williams" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:56.97">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2012-10-14" nation="" />
     <RELAY name="BLU FROG TEAM" nation="USA">
      <CLUB name="BLU FROG TEAM" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ross" nameprefix="" lastname="Bohlken" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lucky" nameprefix="" lastname="Meisenheimer" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marc" nameprefix="" lastname="Middleton" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:19.86">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-11-11" nation="" />
     <RELAY name="RICE AQUATIC MASTERS" nation="USA">
      <CLUB name="RICE AQUATIC MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jay" nameprefix="" lastname="Yarid" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="David" nameprefix="" lastname="Guthrie" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="John" nameprefix="" lastname="Fields" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Bruce" nameprefix="" lastname="Williams" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:50.43">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-12-04" nation="" />
     <RELAY name="VENTURA COUNTY MASTERS" nation="USA">
      <CLUB name="VENTURA COUNTY MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jim" nameprefix="" lastname="McConica" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Glenn" nameprefix="" lastname="Gruber" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Michael" nameprefix="" lastname="Blatt" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Mike" nameprefix="" lastname="Shaffer" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:25.42">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <RELAY name="SWOL 1894" nation="NED">
      <CLUB name="SWOL 1894" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jappie" nameprefix="" lastname="Kuiper" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Mans" nameprefix="" lastname="Buis" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Berkhof" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Harry" nameprefix="" lastname="Dokter" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:39.01">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2017-12-02" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:44.11">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2024-01-06" nation="NED" />
     <RELAY name="SWOL 1894" nation="NED">
      <CLUB name="SWOL 1894" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jappie" nameprefix="" lastname="Kuiper" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Berkhof" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Be" nameprefix="van der" lastname="Ziel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Harry" nameprefix="" lastname="Dokter" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:03.23">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2018-12-02" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Evertjan" nameprefix="" lastname="Masurel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Andr�" nameprefix="" lastname="Pantekoek" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:12:17.60">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:57.97">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Stenungsund" date="2023-03-18" nation="SWE" />
     <RELAY name="G�teborg Sim" nation="SWE">
      <CLUB name="G�teborg Sim" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:16.20">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Firenze" date="2022-03-19" nation="ITA" />
     <RELAY name="DLF Livorno" nation="ITA">
      <CLUB name="DLF Livorno" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:37.70">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Firenze" date="2022-03-20" nation="ITA" />
     <RELAY name="DLF Livorno" nation="ITA">
      <CLUB name="DLF Livorno" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:13.11">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Hodmezovazarvehely" date="2021-09-25" nation="HUN" />
     <RELAY name="T�r�kbalinti senior" nation="HUN">
      <CLUB name="T�r�kbalinti senior" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:58.32">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rapallo" date="2022-04-10" nation="ITA" />
     <RELAY name="Rapallo Nuoto" nation="ITA">
      <CLUB name="Rapallo Nuoto" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:54.44">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-10-11" nation="" />
     <RELAY name="GOLD COAST MASTERS" nation="USA">
      <CLUB name="GOLD COAST MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Keefe" nameprefix="" lastname="Lodwig" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jan" nameprefix="" lastname="Soderstrom" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lee" nameprefix="" lastname="Childs" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="David" nameprefix="" lastname="Quiggin" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:10.51">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-10-22" nation="" />
     <RELAY name="Esporte Cube Pinhei" nation="BRA">
      <CLUB name="Esporte Cube Pinhei" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:19.08">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-11-13" nation="" />
     <RELAY name="Sarasota Sharks" nation="USA">
      <CLUB name="Sarasota Sharks" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:59.48">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-05-25" nation="" />
     <RELAY name="VENTURA COUNTY MASTERS" nation="USA">
      <CLUB name="VENTURA COUNTY MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Steven" nameprefix="" lastname="Heck" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hubie" nameprefix="" lastname="Kerns" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Glenn" nameprefix="" lastname="Gruber" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Bruce" nameprefix="" lastname="Rollins" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:45.48">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-11-06" nation="" />
     <RELAY name="Sarasota Sharks Masters" nation="USA">
      <CLUB name="Sarasota Sharks Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:25.37">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eskilstuna" date="2019-03-23" nation="SWE" />
     <RELAY name="Hellas SK Stockholm" nation="SWE">
      <CLUB name="Hellas SK Stockholm" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:49.33">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Szazhalombatta" date="2020-02-16" nation="HUN" />
     <RELAY name="T�r�kbalinti Senior" nation="HUN">
      <CLUB name="T�r�kbalinti Senior" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:00.26">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2019-10-27" nation="GBR" />
     <RELAY name="Birmingham Masters" nation="GBR">
      <CLUB name="Birmingham Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:57.10">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <RELAY name="Birmingham Masters" nation="GBR">
      <CLUB name="Birmingham Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:14:21.45">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2022-10-28" nation="GBR" />
     <RELAY name="Birmingham Masters" nation="GBR">
      <CLUB name="Birmingham Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:12.76">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-10-08" nation="" />
     <RELAY name="Tamaloais Aquatics Masters" nation="USA">
      <CLUB name="Tamaloais Aquatics Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:37.06">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-10-07" nation="" />
     <RELAY name="Tamalpais Aquatic Masters" nation="USA">
      <CLUB name="Tamalpais Aquatic Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:00.23">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-10-07" nation="" />
     <RELAY name="Tamalpais Aquatic Masters" nation="USA">
      <CLUB name="Tamalpais Aquatic Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:14.65">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-04-02" nation="" />
     <RELAY name="Esporte Clube Pinhei" nation="BRA">
      <CLUB name="Esporte Clube Pinhei" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:11:23.16">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-10-06" nation="" />
     <RELAY name="Tamalpais Aquatic Masters" nation="USA">
      <CLUB name="Tamalpais Aquatic Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:06:54.67">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Palma de Mallorca" date="2017-02-02" nation="ESP" />
     <RELAY name="ESMAS" nation="ESP">
      <CLUB name="ESMAS" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:03:19.42">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2008-02-17" nation="" />
     <RELAY name="JUEI CLUB" nation="JPN">
      <CLUB name="JUEI CLUB" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Isamu" nameprefix="" lastname="Tamura" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hidekazu" nameprefix="" lastname="Tamura" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Hideya" nameprefix="" lastname="Fujii" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Tokushi" nameprefix="" lastname="Komeda" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:15.49">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-05-09" nation="" />
     <RELAY name="NISHINOMIYA SUMIRE" nation="JPN">
      <CLUB name="NISHINOMIYA SUMIRE" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Toshio" nameprefix="" lastname="Yuri" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Takeshi" nameprefix="" lastname="Yasukawa" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Himoru" nameprefix="" lastname="Yoshimoto" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Kazunaga" nameprefix="" lastname="Akutsu" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:52.10">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2014-10-12" nation="" />
     <RELAY name="FLORIDA AQUATIC COMBINED" nation="USA">
      <CLUB name="FLORIDA AQUATIC COMBINED" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rogers" nameprefix="" lastname="Holmes" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="John" nameprefix="" lastname="Corse" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Edwin" nameprefix="" lastname="Graves" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="William" nameprefix="" lastname="Adams" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:21:24.39">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2014-10-10" nation="" />
     <RELAY name="FLORIDA AQUATIC COMBINED" nation="USA">
      <CLUB name="FLORIDA AQUATIC COMBINED" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rogers" nameprefix="" lastname="Holmes" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="William" nameprefix="" lastname="Adams" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Edwin" nameprefix="" lastname="Graves" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="John" nameprefix="" lastname="Corse" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="99" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:40.64">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="Albion WSS (SG)" nation="NED">
      <CLUB name="Albion WSS (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Thomas" nameprefix="" lastname="Verhoeven" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fenna" nameprefix="de" lastname="Groot" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Dinkelberg" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:50.83">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="Albion WSS (SG)" nation="NED">
      <CLUB name="Albion WSS (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Fenna" nameprefix="de" lastname="Groot" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Thomas" nameprefix="" lastname="Verhoeven" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Dinkelberg" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:39.84">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="Albion WSS (SG)" nation="NED">
      <CLUB name="Albion WSS (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Thomas" nameprefix="" lastname="Verhoeven" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fenna" nameprefix="de" lastname="Groot" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Dinkelberg" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:04.06">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="Albion WSS (SG)" nation="NED">
      <CLUB name="Albion WSS (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Fenna" nameprefix="de" lastname="Groot" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Thomas" nameprefix="" lastname="Verhoeven" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Dinkelberg" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:31.48">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <RELAY name="ZVL-1886 Center" nation="NED">
      <CLUB name="ZVL-1886 Center" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Robin" nameprefix="van" lastname="Beek" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Guus" nameprefix="" lastname="Hoogduin" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Karen" nameprefix="" lastname="Stolk" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Silke" nameprefix="" lastname="Molendijk" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:41.34">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2014-01-26" nation="NED" />
     <RELAY name="DWK" nation="NED">
      <CLUB name="DWK" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Nick" nameprefix="van" lastname="Gemert" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marloes" nameprefix="" lastname="Erkens" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Pauline" nameprefix="" lastname="Gouwens" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Merijn" nameprefix="" lastname="Ellenkamp" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:49.19">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="Rotterdam Swimming (SG)" nation="NED">
      <CLUB name="Rotterdam Swimming (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Babette" nameprefix="van der" lastname="Kaaij" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Mark" nameprefix="" lastname="Baars" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Alisha" nameprefix="" lastname="Vieira" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:40.20">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="VZC" nation="NED">
      <CLUB name="VZC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marjolein" nameprefix="" lastname="Delno" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Olaf" nameprefix="" lastname="Achterberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jelle" nameprefix="" lastname="Nap" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Saskia" nameprefix="de" lastname="Jonge" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:05.65">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2014-01-25" nation="NED" />
     <RELAY name="DWK" nation="NED">
      <CLUB name="DWK" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Merijn" nameprefix="" lastname="Ellenkamp" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Nick" nameprefix="van" lastname="Gemert" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Pauline" nameprefix="" lastname="Gouwens" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marion" nameprefix="van den" lastname="Berg" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:16.24">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <RELAY name="DZ&amp;PC" nation="NED">
      <CLUB name="DZ&amp;PC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Am�" nameprefix="" lastname="Hulleman" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Nijholt" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Karin" nameprefix="" lastname="Rijkelijkhuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jelle" nameprefix="" lastname="Betten" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:38.76">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-10-29" nation="GBR" />
     <RELAY name="Bristol Henleaze" nation="GBR">
      <CLUB name="Bristol Henleaze" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:47.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2021-11-22" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novgorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novgorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:40.20">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="VZC" nation="NED">
      <CLUB name="VZC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marjolein" nameprefix="" lastname="Delno" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Olaf" nameprefix="" lastname="Achterberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jelle" nameprefix="" lastname="Nap" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Saskia" nameprefix="de" lastname="Jonge" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:01.17">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2020-11-22" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novograd" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novograd" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:14.19">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Blackpool" date="2022-02-26" nation="GBR" />
     <RELAY name="Trafford Masters" nation="GBR">
      <CLUB name="Trafford Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:38.76">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-10-29" nation="" />
     <RELAY name="Bristol Hen" nation="GBR">
      <CLUB name="Bristol Hen" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:45.63">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-05-21" nation="" />
     <RELAY name="Queendom" nation="JPN">
      <CLUB name="Queendom" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:40.20">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="VZC" nation="NED">
      <CLUB name="VZC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marjolein" nameprefix="" lastname="Delno" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Olaf" nameprefix="" lastname="Achterberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jelle" nameprefix="" lastname="Nap" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Saskia" nameprefix="de" lastname="Jonge" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:01.17">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2020-11-22" nation="" />
     <RELAY name="Tsunami" nation="RUS">
      <CLUB name="Tsunami" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Egor" nameprefix="" lastname="Iogin" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Anton" nameprefix="" lastname="Tishchenko" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Irina" nameprefix="" lastname="Shlemova" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Alina" nameprefix="" lastname="Demkina" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:14.19">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-02-26" nation="" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:44.78">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Nijverdal" date="2013-01-27" nation="NED" />
     <RELAY name="HZ&amp;PC HEERENVEEN" nation="NED">
      <CLUB name="HZ&amp;PC HEERENVEEN" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ren�" nameprefix="" lastname="Beetsma" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Nanda" nameprefix="de" lastname="Vries" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Chantal" nameprefix="" lastname="Nap" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:53.87">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <RELAY name="SwimGym" nation="NED">
      <CLUB name="SwimGym" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Tessa" nameprefix="" lastname="Brouwer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Aleksey" nameprefix="" lastname="Bayevsky" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Andrea" nameprefix="" lastname="Kneppers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="S�bas" nameprefix="van" lastname="Lith" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:45.25">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <RELAY name="SwimGym" nation="NED">
      <CLUB name="SwimGym" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Tessa" nameprefix="" lastname="Brouwer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Aleksey" nameprefix="" lastname="Bayevsky" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Andrea" nameprefix="" lastname="Kneppers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="S�bas" nameprefix="van" lastname="Lith" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:13.05">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Danielle" nameprefix="de" lastname="Boer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Dennis" nameprefix="" lastname="Bos" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fraukje" nameprefix="" lastname="Puts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:38.57">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-24" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Dennis" nameprefix="" lastname="Bos" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Danielle" nameprefix="de" lastname="Boer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fraukje" nameprefix="" lastname="Puts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:37.51">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Saransk" date="2019-11-22" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novgorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novgorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:47.55">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2021-11-17" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novgorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novgorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:36.49">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Getxo" date="2023-06-10" nation="ESP" />
     <RELAY name="Getxo" nation="ESP">
      <CLUB name="Getxo" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:06.82">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Firenze" date="2022-03-19" nation="ITA" />
     <RELAY name="Roma Nuoto Masters" nation="ITA">
      <CLUB name="Roma Nuoto Masters" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:07.91">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2022-10-30" nation="GBR" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:37.51">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-11-22" nation="" />
     <RELAY name="TSUNAMI" nation="RUS">
      <CLUB name="TSUNAMI" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Andrei" nameprefix="" lastname="Kurnosov" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Aleksey" nameprefix="" lastname="Getmanenko" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ekatarina" nameprefix="" lastname="Yudina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Irina" nameprefix="" lastname="Shlemova" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:47.26">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-05-26" nation="" />
     <RELAY name="Wild Rose Swim Club" nation="CAN">
      <CLUB name="Wild Rose Swim Club" nation="CAN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:36.49">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-10-06" nation="" />
     <RELAY name="Getxo" nation="ESP">
      <CLUB name="Getxo" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:56.24">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2013-11-24" nation="" />
     <RELAY name="PHOENIX SWIM CLUB" nation="USA">
      <CLUB name="PHOENIX SWIM CLUB" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Noriko" nameprefix="" lastname="Inada" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jeff" nameprefix="" lastname="Commings" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erin" nameprefix="" lastname="Campbell" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jan" nameprefix="" lastname="Konarzewski" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:07.91">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-10-30" nation="" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:46.71">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-27" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jeroen" nameprefix="" lastname="Zelsmann" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:57.61">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Rotterdam" date="2020-01-26" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Joan" nameprefix="" lastname="Kentrop" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:58.63">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Danielle" nameprefix="de" lastname="Boer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:20.45">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Terneuzen" date="2018-01-21" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:53.25">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-19" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fraukje" nameprefix="" lastname="Puts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:40.86">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="St. Petersburg" date="2015-11-28" nation="RUS" />
     <RELAY name="Neva Stars" nation="RUS">
      <CLUB name="Neva Stars" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:50.35">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2021-11-14" nation="RUS" />
     <RELAY name="Mad Wave" nation="RUS">
      <CLUB name="Mad Wave" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:48.27">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2017-10-27" nation="GBR" />
     <RELAY name="Basingstoke Masters" nation="GBR">
      <CLUB name="Basingstoke Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:10.95">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Roma" date="2018-04-21" nation="ITA" />
     <RELAY name="Brescia aquare Mafeco" nation="ITA">
      <CLUB name="Brescia aquare Mafeco" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:19.38">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Ostia" date="2023-03-12" nation="ITA" />
     <RELAY name="Circolo Canottieri Aniene" nation="ITA">
      <CLUB name="Circolo Canottieri Aniene" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:40.07">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-11-11" nation="" />
     <RELAY name="Tsunami" nation="RUS">
      <CLUB name="Tsunami" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Andrey" nameprefix="" lastname="Kurnosov" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:50.35">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-11-14" nation="" />
     <RELAY name="Mad Wave" nation="RUS">
      <CLUB name="Mad Wave" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:46.01">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2009-11-21" nation="" />
     <RELAY name="COLORADO MASTERS" nation="USA">
      <CLUB name="COLORADO MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chris" nameprefix="" lastname="O'sullivan" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Sheri" nameprefix="" lastname="Hart" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:05.01">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-05-07" nation="" />
     <RELAY name="JSS Fukai" nation="JPN">
      <CLUB name="JSS Fukai" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:19.38">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-03-12" nation="" />
     <RELAY name="CC Aniene" nation="ITA">
      <CLUB name="CC Aniene" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:51.85">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Oss" date="2022-09-25" nation="NED" />
     <RELAY name="Zpc Amersfoort" nation="NED">
      <CLUB name="Zpc Amersfoort" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jeroen" nameprefix="" lastname="Zelsmann" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:05.42">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Zwolle" date="2019-01-26" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:10.79">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Nijverdal" date="2013-01-27" nation="NED" />
     <RELAY name="AZ&amp;PC" nation="NED">
      <CLUB name="AZ&amp;PC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ron" nameprefix="" lastname="Korzelius" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:31.75">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2014-06-28" nation="NED" />
     <RELAY name="AZ&amp;PC" nation="NED">
      <CLUB name="AZ&amp;PC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Stefan" nameprefix="" lastname="Dortmond" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:13.45">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Nijverdal" date="2013-01-25" nation="NED" />
     <RELAY name="AZ&amp;PC" nation="NED">
      <CLUB name="AZ&amp;PC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ron" nameprefix="" lastname="Korzelius" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:46.08">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2016-10-28" nation="GBR" />
     <RELAY name="East Leeds" nation="GBR">
      <CLUB name="East Leeds" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:58.12">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2023-10-28" nation="GBR" />
     <RELAY name="Woking" nation="GBR">
      <CLUB name="Woking" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:57.51">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2021-10-30" nation="GBR" />
     <RELAY name="East Leeds" nation="GBE">
      <CLUB name="East Leeds" nation="GBE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:25.65">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2022-10-28" nation="GBR" />
     <RELAY name="Woking" nation="GBR">
      <CLUB name="Woking" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:54.52">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Pomezia" date="2023-01-29" nation="ITA" />
     <RELAY name="Circolo Canottieri Aniene" nation="ITA">
      <CLUB name="Circolo Canottieri Aniene" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:45.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-04-16" nation="" />
     <RELAY name="Edge" nation="JPN">
      <CLUB name="Edge" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:55.87">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-04-16" nation="" />
     <RELAY name="Edge" nation="JPN">
      <CLUB name="Edge" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:56.10">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2014-12-14" nation="" />
     <RELAY name="NORTH CAROLINA MASTERS" nation="USA">
      <CLUB name="NORTH CAROLINA MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Henry" nameprefix="" lastname="Stewart" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Sue" nameprefix="" lastname="Walsh" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jonathan" nameprefix="" lastname="Klein" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:19.84">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-03-18" nation="" />
     <RELAY name="North Carolina Masters" nation="USA">
      <CLUB name="North Carolina Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:36.91">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-10-11" nation="" />
     <RELAY name="ILLINOIS MASTERS" nation="USA">
      <CLUB name="ILLINOIS MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Liz" nameprefix="" lastname="Dillmann" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="David" nameprefix="" lastname="Sims" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Andrea" nameprefix="" lastname="Block" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jim" nameprefix="" lastname="Tuchler" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:53.75">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:10.06">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:13.40">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:48.46">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:25.75">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:53.75">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:08.89">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Brescia" date="2023-01-29" nation="ITA" />
     <RELAY name="Acqua1 Village SSD" nation="ITA">
      <CLUB name="Acqua1 Village SSD" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:13.40">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:48.46">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Heerenveen" date="2023-02-18" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:25.75">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:52.68">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-11-14" nation="" />
     <RELAY name="NORTH TEXAS LONESTARS" nation="USA">
      <CLUB name="NORTH TEXAS LONESTARS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Doug" nameprefix="" lastname="Martin" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Tom" nameprefix="" lastname="Barton" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Christina" nameprefix="" lastname="Mckelvey" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lynn" nameprefix="" lastname="Morrison" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:04.82">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-07-12" nation="" />
     <RELAY name="NOVAQUATICS MASTERS" nation="USA">
      <CLUB name="NOVAQUATICS MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jamie" nameprefix="" lastname="Fowler" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Henry" nameprefix="" lastname="Vehovec" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Katie" nameprefix="" lastname="Osborne" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Veronica" nameprefix="" lastname="Hibben" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:13.40">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-19" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:43.20">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-12-13" nation="" />
     <RELAY name="OREGON MASTERS" nation="USA">
      <CLUB name="OREGON MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Karen" nameprefix="" lastname="Andrus-Hughes" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Colette" nameprefix="" lastname="Crabbe" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Allen" nameprefix="" lastname="Stark" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:25.75">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2023-02-17" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:15.40">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Rotterdam" date="2020-01-25" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:38.89">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Steenwijk" date="2019-09-14" nation="NED" />
     <RELAY name="Psv" nation="NED">
      <CLUB name="Psv" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Evertjan" nameprefix="" lastname="Masurel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:18.73">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:54.71">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2014-12-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:12:07.16">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Heerenveen" date="2015-01-23" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:12.77">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:32.69">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Lodi" date="2023-02-12" nation="ITA" />
     <RELAY name="Aly sport ASD" nation="ITA">
      <CLUB name="Aly sport ASD" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:18.73">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Terneuzen" date="2018-01-20" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:47.93">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2023-10-29" nation="GBR" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:11:47.24">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Bordeaux" date="2022-01-30" nation="FRA" />
     <RELAY name="Bordeaux ETU club" nation="FRA">
      <CLUB name="Bordeaux ETU club" nation="FRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:07.33">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-10-09" nation="" />
     <RELAY name="Tamalpais Masters" nation="USA">
      <CLUB name="Tamalpais Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:22.04">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-09-27" nation="" />
     <RELAY name="TAMALPAIS AQUATIC MASTERS" nation="USA">
      <CLUB name="TAMALPAIS AQUATIC MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kenneth" nameprefix="" lastname="Frost" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nancy" nameprefix="" lastname="Ridout" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:40.10">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-10-08" nation="" />
     <RELAY name="Tamalpais Masters" nation="USA">
      <CLUB name="Tamalpais Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:21.37">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-10-11" nation="" />
     <RELAY name="TAMALPAIS AQUATIC MASTERS" nation="USA">
      <CLUB name="TAMALPAIS AQUATIC MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kenneth" nameprefix="" lastname="Frost" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nancy" nameprefix="" lastname="Ridout" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:54.11">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-09-27" nation="" />
     <RELAY name="TAMALPAIS AQUATIC MASTERS" nation="USA">
      <CLUB name="TAMALPAIS AQUATIC MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kenneth" nameprefix="" lastname="Frost" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Nancy" nameprefix="" lastname="Ridout" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:03:06.81">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Funchal" date="2023-11-19" nation="POR" />
     <RELAY name="Psv" nation="NED">
      <CLUB name="Psv" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:07.47">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Veldhoven" date="2015-02-08" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:37.53">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2012-03-17" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Aloys" nameprefix="" lastname="Geurts" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Cor" nameprefix="" lastname="Sprengers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:29.92">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2023-11-26" nation="NED" />
     <RELAY name="Psv" nation="NED">
      <CLUB name="Psv" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Gonnie" nameprefix="" lastname="Bak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Henk" nameprefix="" lastname="Maessen" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:14:49.10">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-12-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jan" nameprefix="" lastname="Nuijten" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:43.90">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <RELAY name="Birmingham Masters" nation="GBR">
      <CLUB name="Birmingham Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:00.58">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Aartselaar" date="2016-05-21" nation="BEL" />
     <RELAY name="AZSC" nation="BEL">
      <CLUB name="AZSC" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:19.86">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2022-10-29" nation="GBR" />
     <RELAY name="Birmingham Masters" nation="GBR">
      <CLUB name="Birmingham Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:12.41">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Maastricht" date="2017-01-22" nation="NED" />
     <RELAY name="Antwerpse Zwemclub Scaldis" nation="BEL">
      <CLUB name="Antwerpse Zwemclub Scaldis" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jozef" nameprefix="van" lastname="Roy" gender="M" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Joseph" nameprefix="" lastname="Meyten" gender="M" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Eliane" nameprefix="" lastname="Pellis" gender="F" nation="BEL" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:14:26.47">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2022-10-30" nation="GBR" />
     <RELAY name="Birmingham Masters" nation="GBR">
      <CLUB name="Birmingham Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:26.62">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-01-27" nation="" />
     <RELAY name="ST. KANSAI" nation="JPN">
      <CLUB name="ST. KANSAI" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Fusako" nameprefix="" lastname="Hirooka" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Yoshiko" nameprefix="" lastname="Osaki" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Chitoshi" nameprefix="" lastname="Konishi" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Yoshiyuki" nameprefix="" lastname="Funahashi" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:57.97">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-10-03" nation="" />
     <RELAY name="OREGON MASTERS" nation="USA">
      <CLUB name="OREGON MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Janet" nameprefix="" lastname="Gettling" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Margaret" nameprefix="" lastname="Toppel" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:00.74">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-11-12" nation="" />
     <RELAY name="OREGON MASTERS" nation="USA">
      <CLUB name="OREGON MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Joy" nameprefix="" lastname="Ward" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Margaret" nameprefix="" lastname="Toppel" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:59.56">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-11-11" nation="" />
     <RELAY name="OREGON MASTERS" nation="USA">
      <CLUB name="OREGON MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Janet" nameprefix="" lastname="Gettling" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Joy" nameprefix="" lastname="Ward" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:14:26.47">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-10-30" nation="" />
     <RELAY name="Birmingham Masters" nation="GBR">
      <CLUB name="Birmingham Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="SCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:03:32.71">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2018-02-11" nation="" />
     <RELAY name="SUNWAY YOKOHAMA" nation="JPN">
      <CLUB name="SUNWAY YOKOHAMA" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Meiko" nameprefix="" lastname="Kamashita" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kaizo" nameprefix="" lastname="Watanabe" gender="X" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Minoru" nameprefix="" lastname="Nagashima" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:02.42">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-04-22" nation="" />
     <RELAY name="Warringah Masters" nation="AUS">
      <CLUB name="Warringah Masters" nation="AUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:05.56">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-10-21" nation="" />
     <RELAY name="SUNWAY YOKOHAMA" nation="JPN">
      <CLUB name="SUNWAY YOKOHAMA" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Meiko" nameprefix="" lastname="Kamashita" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kaizo" nameprefix="" lastname="Watanabe" gender="X" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Shigeko" nameprefix="" lastname="Tanaka" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Minoru" nameprefix="" lastname="Nagashima" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:38.12">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-05-31" nation="" />
     <RELAY name="SAPPORO MST" nation="JPN">
      <CLUB name="SAPPORO MST" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Fumi" nameprefix="" lastname="Murata" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Naka" nameprefix="" lastname="Fukuoka" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Toshikazu" nameprefix="" lastname="Tateda" gender="X" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Yoshiro" nameprefix="" lastname="Obata" gender="X" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:23:00.65">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2016-12-17" nation="" />
     <RELAY name="FLORIDA AQUATIC COMBINED" nation="USA">
      <CLUB name="FLORIDA AQUATIC COMBINED" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Edwin" nameprefix="" lastname="Graves" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="John" nameprefix="" lastname="Corse" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Joan" nameprefix="" lastname="Campbell" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Betty" nameprefix="" lastname="Lorenzi" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="99" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:51.98">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-03" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kimberley" nameprefix="" lastname="Albers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Isabelle" nameprefix="" lastname="Massar" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Manon" nameprefix="van" lastname="Strien" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Anja" nameprefix="van der" lastname="Hout" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:05.15">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="Hieronymus" nation="NED">
      <CLUB name="Hieronymus" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Valesca" nameprefix="van den" lastname="Bogert" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Selene" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Christel" nameprefix="" lastname="Brugmans" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nadja" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:06.67">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <RELAY name="Hieronymus" nation="NED">
      <CLUB name="Hieronymus" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marlijn" nameprefix="" lastname="Hendriksen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Eva" nameprefix="van" lastname="Ginneken" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Nadja" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Selene" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:36.61">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="Hieronymus" nation="NED">
      <CLUB name="Hieronymus" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Nadja" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Valesca" nameprefix="van den" lastname="Bogert" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Selene" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Roos" nameprefix="" lastname="Englebert" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:07.56">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <RELAY name="Hieronymus" nation="NED">
      <CLUB name="Hieronymus" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Selene" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Nadja" nameprefix="" lastname="Wortel" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Valesca" nameprefix="van den" lastname="Bogert" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Roos" nameprefix="" lastname="Englebert" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:51.61">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Londen" date="2016-05-26" nation="GBR" />
     <RELAY name="De Dinkel" nation="NED">
      <CLUB name="De Dinkel" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Karin" nameprefix="" lastname="Hidding" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Anique" nameprefix="" lastname="Willeme" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Silke" nameprefix="" lastname="Oude Weernink" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marlies" nameprefix="" lastname="Reinders" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:04.09">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Londen" date="2016-05-27" nation="GBR" />
     <RELAY name="De Dinkel" nation="NED">
      <CLUB name="De Dinkel" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Silke" nameprefix="" lastname="Oude Weernink" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Karin" nameprefix="" lastname="Hidding" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anique" nameprefix="" lastname="Willeme" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marlies" nameprefix="" lastname="Reinders" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:06.21">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Manon" nameprefix="van" lastname="Strien" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Isabelle" nameprefix="" lastname="Massar" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:39.75">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2017-05-07" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Manon" nameprefix="van" lastname="Strien" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Nicole" nameprefix="" lastname="Bennis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Isabelle" nameprefix="" lastname="Massar" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:25.00">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Nicole" nameprefix="" lastname="Bennis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Manon" nameprefix="van" lastname="Strien" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Isabelle" nameprefix="" lastname="Massar" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:50.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Kazan" date="2015-08-14" nation="RUS" />
     <RELAY name="NEVA STARS" nation="RUS">
      <CLUB name="NEVA STARS" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Evgenia" nameprefix="" lastname="Karetina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ekaterina" nameprefix="" lastname="Shershen" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anna" nameprefix="" lastname="Kuzmicheva" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Anna" nameprefix="" lastname="Polyakova" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:00.05">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Kazan" date="2015-08-14" nation="RUS" />
     <RELAY name="NEVA STARS" nation="RUS">
      <CLUB name="NEVA STARS" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Evgenia" nameprefix="" lastname="Karetina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Anna" nameprefix="" lastname="Kuzmicheva" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anna" nameprefix="" lastname="Polyakova" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ekaterina" nameprefix="" lastname="Shershen" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:03.63">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-04" nation="GBR" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:42.20">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="St. Petersburg" date="2022-02-24" nation="RUS" />
     <RELAY name="Tsunami Nizhniy" nation="RUS">
      <CLUB name="Tsunami Nizhniy" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:02.70">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Braunschweig" date="2016-02-27" nation="GER" />
     <RELAY name="SG Dortmund" nation="GER">
      <CLUB name="SG Dortmund" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kerstin" nameprefix="" lastname="Lange" gender="F" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Mandy" nameprefix="" lastname="Blum" gender="F" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrina" nameprefix="" lastname="Miede" gender="F" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jennifer" nameprefix="" lastname="Thater" gender="F" nation="GER" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:50.28">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2016-10-16" nation="" />
     <RELAY name="CMC SC" nation="JPN">
      <CLUB name="CMC SC" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Natsuki" nameprefix="" lastname="Hasegawa" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Natsumi" nameprefix="" lastname="Mizuochi" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Sanae" nameprefix="" lastname="Nawata" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ayaka" nameprefix="" lastname="Kawabata" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:00.05">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-08-14" nation="" />
     <RELAY name="NEVA STARS" nation="RUS">
      <CLUB name="NEVA STARS" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Evgenia" nameprefix="" lastname="Karetina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Anna" nameprefix="" lastname="Kuzmicheva" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anna" nameprefix="" lastname="Polyakova" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ekaterina" nameprefix="" lastname="Shershen" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:00.96">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-12-11" nation="" />
     <RELAY name="Linx racing Team" nation="JPN">
      <CLUB name="Linx racing Team" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:30.81">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-12-11" nation="" />
     <RELAY name="Linx Racing Team" nation="JPN">
      <CLUB name="Linx Racing Team" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:58.97">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-12-12" nation="" />
     <RELAY name="Linx Racing Team" nation="JPN">
      <CLUB name="Linx Racing Team" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:54.76">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Nicole" nameprefix="" lastname="Bennis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lauren" nameprefix="van" lastname="IJll" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lisa" nameprefix="" lastname="Klatten" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:06.24">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lauren" nameprefix="van" lastname="IJll" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Nicole" nameprefix="" lastname="Bennis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lisa" nameprefix="" lastname="Klatten" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:07.52">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Nicole" nameprefix="" lastname="Bennis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Mabel" nameprefix="" lastname="Sulic" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:39.05">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Mabel" nameprefix="" lastname="Sulic" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Nicole" nameprefix="" lastname="Bennis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Leonie" nameprefix="van" lastname="Noort" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:32.87">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-02" nation="NED" />
     <RELAY name="Het Y" nation="NED">
      <CLUB name="Het Y" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Bravo" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Cynthia" nameprefix="" lastname="Noordermeer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ana-Lara" nameprefix="da" lastname="Silva" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Evelien" nameprefix="" lastname="Sohl" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:49.03">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Kazan" date="2015-08-14" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novosibirsk" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novosibirsk" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Svetlana" nameprefix="" lastname="Kniaginina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Alla" nameprefix="" lastname="Feoktistova" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Liubov" nameprefix="" lastname="Yudina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Irina" nameprefix="" lastname="Shlemova" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:03.78">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="No Stars Swim Club" nation="UKR">
      <CLUB name="No Stars Swim Club" nation="UKR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:04.10">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Swansea" date="2019-06-15" nation="GBR" />
     <RELAY name="Birmingham Masters" nation="GBR">
      <CLUB name="Birmingham Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:35.76">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Magdeburg" date="2017-06-17" nation="GER" />
     <RELAY name="Berliner TSC" nation="GER">
      <CLUB name="Berliner TSC" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:11.39">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Swansea" date="2019-06-15" nation="GBR" />
     <RELAY name="Birmingham Masters" nation="GBR">
      <CLUB name="Birmingham Masters" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:49.03">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-08-14" nation="" />
     <RELAY name="TSUNAMI" nation="RUS">
      <CLUB name="TSUNAMI" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Svetlana" nameprefix="" lastname="Kniaginina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Alla" nameprefix="" lastname="Feoktistova" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Liubov" nameprefix="" lastname="Yudina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Irina" nameprefix="" lastname="Shlemova" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:59.41">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-08-09" nation="" />
     <RELAY name="Team Go Mai Way" nation="JPN">
      <CLUB name="Team Go Mai Way" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:04.10">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-06-15" nation="" />
     <RELAY name="BIRMINGHAM MASTERS" nation="GBR">
      <CLUB name="BIRMINGHAM MASTERS" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Katie" nameprefix="" lastname="Walker-stabeler" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Lane" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anna" nameprefix="" lastname="Mccall" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Justine" nameprefix="" lastname="Clark" gender="F" nation="GBR" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:35.76">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-06-17" nation="" />
     <RELAY name="BERLINER TSC" nation="GER">
      <CLUB name="BERLINER TSC" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Andrea" nameprefix="" lastname="Kutz" gender="F" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Kutz" gender="F" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Nadine" nameprefix="" lastname="Stresing" gender="F" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Josephine" nameprefix="" lastname="Dunger" gender="F" nation="GER" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:10.37">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-11-02" nation="" />
     <RELAY name="Potiguar TNT Masters" nation="BRA">
      <CLUB name="Potiguar TNT Masters" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:54.42">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2004-02-15" nation="NED" />
     <RELAY name="AZ&amp;PC" nation="NED">
      <CLUB name="AZ&amp;PC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marja" nameprefix="" lastname="Bloemzaad" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Petra" nameprefix="" lastname="Casteleijn-Frowijn" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:11.62">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Kranj" date="2018-09-02" nation="SLO" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:23.88">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:52.88">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:53.86">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-05" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marije" nameprefix="van" lastname="Manen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:51.91">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Tsunami Nizhniy" nation="RUS">
      <CLUB name="Tsunami Nizhniy" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:06.57">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Gera" date="2016-04-15" nation="GER" />
     <RELAY name="Berliner TSC" nation="GER">
      <CLUB name="Berliner TSC" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Oxana" nameprefix="" lastname="Bronitskaia" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marta" nameprefix="" lastname="Rumyantseva" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ekatarina" nameprefix="" lastname="Yudina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Liubov" nameprefix="" lastname="Yudina" gender="F" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:12.31">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-04" nation="GBR" />
     <RELAY name="Basingstoke" nation="GBR">
      <CLUB name="Basingstoke" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:52.88">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:17.25">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <RELAY name="Basingstoke" nation="GBR">
      <CLUB name="Basingstoke" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:48.44">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2006-08-08" nation="" />
     <RELAY name="TEAM TYR" nation="USA">
      <CLUB name="TEAM TYR" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Sheri" nameprefix="" lastname="Hart" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Collette" nameprefix="" lastname="Sappey" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anna" nameprefix="" lastname="Pettis-Scott" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Susan" nameprefix="von der" lastname="Lippe" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:02.92">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-08-04" nation="" />
     <RELAY name="North Carolina Masters" nation="USA">
      <CLUB name="North Carolina Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:06.90">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-06-14" nation="" />
     <RELAY name="NORTH CAROLINA MASTERS" nation="USA">
      <CLUB name="NORTH CAROLINA MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Erika" nameprefix="" lastname="Braun" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jen" nameprefix="" lastname="Stringer" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Alicia" nameprefix="" lastname="Uhl" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Kerry" nameprefix="" lastname="Lindauer" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:40.42">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-08-20" nation="" />
     <RELAY name="North Carolina Masters" nation="USA">
      <CLUB name="North Carolina Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:17.25">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-06-03" nation="" />
     <RELAY name="Basingstoke" nation="GBR">
      <CLUB name="Basingstoke" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:58.66">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Barbara" nameprefix="van" lastname="Rhijn" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jenny" nameprefix="" lastname="Bergwerff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:15.91">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jeanne" nameprefix="" lastname="Petit" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:25.78">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:58.55">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Gudule" nameprefix="van der" lastname="Meer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Trudy" nameprefix="" lastname="Ketting-Klaassen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jeanne" nameprefix="" lastname="Petit" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:42.63">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kirsten" nameprefix="" lastname="Cameron" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Katrin" nameprefix="" lastname="Pennings" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Liselotte" nameprefix="" lastname="Joling" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Carla" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:58.66">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Barbara" nameprefix="van" lastname="Rhijn" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jenny" nameprefix="" lastname="Bergwerff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:11.41">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="masters soerlandet" nation="NOR">
      <CLUB name="masters soerlandet" nation="NOR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:25.78">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lidia" nameprefix="van" lastname="Bon-Rosenbrand" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:54.41">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Kristiansand" date="2020-01-25" nation="NOR" />
     <RELAY name="Sorlandet Masters" nation="NOR">
      <CLUB name="Sorlandet Masters" nation="NOR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:08.34">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <RELAY name="Harrogate &amp; District SC" nation="GBR">
      <CLUB name="Harrogate &amp; District SC" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:54.10">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-08-05" nation="" />
     <RELAY name="North Carolina Masters" nation="USA">
      <CLUB name="North Carolina Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:08.87">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-08-04" nation="" />
     <RELAY name="Club Tribe" nation="USA">
      <CLUB name="Club Tribe" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:20.68">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2013-03-14" nation="" />
     <RELAY name="CAPE TOWN MASTERS" nation="RSA">
      <CLUB name="CAPE TOWN MASTERS" nation="RSA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Sanderina" nameprefix="" lastname="Kruger" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Cecilia" nameprefix="" lastname="Stanford" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Edith" nameprefix="" lastname="Ottermann" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Perry-Ann" nameprefix="" lastname="Cadiz" gender="F" nation="RSA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:54.41">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2020-01-25" nation="" />
     <RELAY name="MASTERS SORLANDET" nation="NOR">
      <CLUB name="MASTERS SORLANDET" nation="NOR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lise" nameprefix="" lastname="Lothe" gender="F" nation="NOR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Anette" nameprefix="" lastname="Soerensen" gender="F" nation="NOR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Janne" nameprefix="" lastname="Thorstensen" gender="F" nation="NOR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Fuglestveit" gender="F" nation="NOR" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:34.53">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-07-07" nation="" />
     <RELAY name="CONEJO VALLEY MASTERS" nation="USA">
      <CLUB name="CONEJO VALLEY MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jill" nameprefix="" lastname="Gellatly" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Becky" nameprefix="" lastname="Cleavenger" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Eve" nameprefix="" lastname="Maidenberg" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Leslie" nameprefix="" lastname="Daland-james" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:13.23">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-08" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:36.22">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Katrin" nameprefix="" lastname="Pennings" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Katja" nameprefix="de" lastname="Beer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:00.73">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Saskia" nameprefix="" lastname="Phaff" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:04.52">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Krupiarz" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:11:18.86">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:11.09">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Kranj" date="2018-09-05" nation="SLO" />
     <RELAY name="Danderyds Sim Club" nation="SWE">
      <CLUB name="Danderyds Sim Club" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Asa" nameprefix="" lastname="Inde" gender="F" nation="SWE" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:26.23">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <RELAY name="Cercle De Natation Sportcity Woluwe" nation="BEL">
      <CLUB name="Cercle De Natation Sportcity Woluwe" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Pierrette" nameprefix="" lastname="Michel" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Colette" nameprefix="" lastname="Crabb�" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Claire" nameprefix="" lastname="Anthony" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nathalie" nameprefix="" lastname="Blondeel" gender="F" nation="BEL" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:57.76">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <RELAY name="Cercle De Natation Sportcity Woluwe" nation="BEL">
      <CLUB name="Cercle De Natation Sportcity Woluwe" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Colette" nameprefix="" lastname="Crabb�" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Pierrette" nameprefix="" lastname="Michel" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Claire" nameprefix="" lastname="Anthony" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nathalie" nameprefix="" lastname="Blondeel" gender="F" nation="BEL" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:34.98">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="Cercle De Natation Sportcity Woluwe" nation="BEL">
      <CLUB name="Cercle De Natation Sportcity Woluwe" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Pierrette" nameprefix="" lastname="Michel" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Colette" nameprefix="" lastname="Crabb�" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Claire" nameprefix="" lastname="Anthony" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nathalie" nameprefix="" lastname="Blondeel" gender="F" nation="BEL" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:52.10">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <RELAY name="Gateshead &amp; Wickham" nation="GBR">
      <CLUB name="Gateshead &amp; Wickham" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:00.75">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2018-03-17" nation="" />
     <RELAY name="CAPE TOWN MASTERS" nation="RSA">
      <CLUB name="CAPE TOWN MASTERS" nation="RSA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Edith" nameprefix="" lastname="Ottermann" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Sanderina" nameprefix="" lastname="Kruger" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Diane" nameprefix="" lastname="Coetzee" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Cecilia" nameprefix="" lastname="Stanford" gender="F" nation="RSA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:19.90">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-03-16" nation="" />
     <RELAY name="CAPE TOWN MASTERS" nation="RSA">
      <CLUB name="CAPE TOWN MASTERS" nation="RSA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Diane" nameprefix="" lastname="Coetzee" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Cecilia" nameprefix="" lastname="Stanford" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Edith" nameprefix="" lastname="Ottermann" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Sanderina" nameprefix="" lastname="Kruger" gender="F" nation="RSA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:36.74">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-07-21" nation="" />
     <RELAY name="NORTH TEXAS LONESTAR" nation="USA">
      <CLUB name="NORTH TEXAS LONESTAR" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Stephanie" nameprefix="" lastname="Stone" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kristin" nameprefix="" lastname="Henderson" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lynn" nameprefix="" lastname="Morrison" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jeannie" nameprefix="" lastname="Woolslayer" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:19.05">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-02-27" nation="" />
     <RELAY name="CAPE TOWN MASTERS" nation="RSA">
      <CLUB name="CAPE TOWN MASTERS" nation="RSA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Diane" nameprefix="" lastname="Coetzee" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Gail" nameprefix="" lastname="Mccarney" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Cecilia" nameprefix="" lastname="Stanford" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Sanderina" nameprefix="" lastname="Kruger" gender="F" nation="RSA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:13.61">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2016-02-21" nation="" />
     <RELAY name="CAPE TOWN MASTERS" nation="RSA">
      <CLUB name="CAPE TOWN MASTERS" nation="RSA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Cecilia" nameprefix="" lastname="Stanford" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Gail" nameprefix="" lastname="Mccarney" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Diane" nameprefix="" lastname="Coetzee" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Sanderina" nameprefix="" lastname="Kruger" gender="F" nation="RSA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:30.19">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Krupiarz" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:05.98">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2013-09-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Krupiarz" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:39.58">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:43.79">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Krupiarz" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:12:25.08">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:29.53">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="NeuK�lln Berlin" nation="GER">
      <CLUB name="NeuK�lln Berlin" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:47.19">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="London" date="2016-05-29" nation="GBR" />
     <RELAY name="Spencer Swim Team" nation="GBR">
      <CLUB name="Spencer Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Janet" nameprefix="" lastname="Brown" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Diane" nameprefix="" lastname="Ford" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Amanda" nameprefix="" lastname="Heath" gender="F" nation="GBR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jean" nameprefix="" lastname="Howard Jones" gender="F" nation="GBR" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:39.58">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:17.26">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Aberdeen" date="2022-06-19" nation="GBR" />
     <RELAY name="Spencer Swim Team" nation="GBR">
      <CLUB name="Spencer Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:12:25.08">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:14.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-01-20" nation="USA" />
     <RELAY name="Lone Star Masters" nation="USA">
      <CLUB name="Lone Star Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:34.78">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-01-20" nation="USA" />
     <RELAY name="Lone Star Masters" nation="USA">
      <CLUB name="Lone Star Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:26.29">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-06-12" nation="" />
     <RELAY name="Sarasota Sharks" nation="USA">
      <CLUB name="Sarasota Sharks" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:17.26">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-06-19" nation="" />
     <RELAY name="Spencer" nation="GBR">
      <CLUB name="Spencer" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:12:25.08">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ineke" nameprefix="" lastname="Weekers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Esther" nameprefix="van" lastname="Lohuizen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:03:47.00">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Carla" nameprefix="" lastname="Hensen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Gonnie" nameprefix="" lastname="Bak" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:10.84">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Carla" nameprefix="" lastname="Hensen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:50.07">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-07" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Annie" nameprefix="" lastname="Smits" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:22.93">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Liesbeth" nameprefix="ter" lastname="Laak-Braun" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:18:39.49">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:03:10.24">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Kranj" date="2007-08-29" nation="SLO" />
     <RELAY name="SOIK HELLAS" nation="SWE">
      <CLUB name="SOIK HELLAS" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:36.21">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Riccione" date="2012-06-14" nation="ITA" />
     <RELAY name="SIMKLUBBEN NAUTILUS" nation="SWE">
      <CLUB name="SIMKLUBBEN NAUTILUS" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kerstin" nameprefix="" lastname="Gj�res" gender="F" nation="SWE" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Britt" nameprefix="" lastname="Grilli" gender="F" nation="SWE" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Harriet" nameprefix="" lastname="Bure" gender="F" nation="SWE" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Eva-Britt" nameprefix="" lastname="Widahl" gender="F" nation="SWE" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:00.29">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Swansea" date="2019-06-15" nation="GBR" />
     <RELAY name="Spencer Swim Team" nation="GBR">
      <CLUB name="Spencer Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:21.15">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Swansea" date="2019-06-16" nation="GBR" />
     <RELAY name="Spencer Swim Team" nation="GBR">
      <CLUB name="Spencer Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:18:39.49">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:52.72">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-06-05" nation="" />
     <RELAY name="St Kansai" nation="JPN">
      <CLUB name="St Kansai" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:23.94">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-06-04" nation="" />
     <RELAY name="St Kansai" nation="JPN">
      <CLUB name="St Kansai" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:36.85">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-07-31" nation="" />
     <RELAY name="St. Kansai" nation="JPN">
      <CLUB name="St. Kansai" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:52.67">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-06-18" nation="" />
     <RELAY name="Miami Masters" nation="USA">
      <CLUB name="Miami Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:15:05.19">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-11-27" nation="" />
     <RELAY name="Miami Masters" nation="USA">
      <CLUB name="Miami Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="F" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:05:47.05">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-02-22" nation="" />
     <RELAY name="SUKOYAKA ST" nation="JPN">
      <CLUB name="SUKOYAKA ST" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Masako" nameprefix="" lastname="Kusume" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Masako" nameprefix="" lastname="Otsuka" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Toshiko" nameprefix="" lastname="Amano" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Chiyoko" nameprefix="" lastname="Takizawa" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:53.02">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-08-05" nation="" />
     <RELAY name="SAPPORO MASTERS" nation="JPN">
      <CLUB name="SAPPORO MASTERS" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Sumiko" nameprefix="" lastname="Kuji" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Naka" nameprefix="" lastname="Fukuoka" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Haruko" nameprefix="" lastname="Sasaki" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fumi" nameprefix="" lastname="Murata" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="99" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:37.66">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-07" nation="NED" />
     <RELAY name="Albion d&apos;ELFT (SG)" nation="NED">
      <CLUB name="Albion d&apos;ELFT (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:50.26">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <RELAY name="Albion d&apos;ELFT (SG)" nation="NED">
      <CLUB name="Albion d&apos;ELFT (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jordi" nameprefix="van der" lastname="Weel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:45.69">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-05-05" nation="NED" />
     <RELAY name="LZ 1886" nation="NED">
      <CLUB name="LZ 1886" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lars" nameprefix="" lastname="Sieval" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kristiaan" nameprefix="" lastname="Lenos" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Joost" nameprefix="" lastname="Rijntjes" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Sjoerd" nameprefix="" lastname="Sieval" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:11.22">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2013-05-04" nation="NED" />
     <RELAY name="Octopus" nation="NED">
      <CLUB name="Octopus" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Albert" nameprefix="van" lastname="Piekeren" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Roald" nameprefix="" lastname="Blok" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Emile" nameprefix="" lastname="Manni" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Floris" nameprefix="" lastname="Manni" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:39.26">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-05-03" nation="NED" />
     <RELAY name="LZ 1886" nation="NED">
      <CLUB name="LZ 1886" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lars" nameprefix="" lastname="Sieval" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Joost" nameprefix="" lastname="Rijntjes" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Sjoerd" nameprefix="" lastname="Sieval" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Kristiaan" nameprefix="" lastname="Lenos" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:38.74">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <RELAY name="Feijenoord Albion Zwemclub" nation="NED">
      <CLUB name="Feijenoord Albion Zwemclub" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jordi" nameprefix="van der" lastname="Weel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:50.00">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <RELAY name="Feijenoord Albion Zwemclub" nation="NED">
      <CLUB name="Feijenoord Albion Zwemclub" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jordi" nameprefix="van der" lastname="Weel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:37.83">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <RELAY name="Albion d&apos;ELFT (SG)" nation="NED">
      <CLUB name="Albion d&apos;ELFT (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:02.05">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <RELAY name="Feijenoord Albion Zwemclub" nation="NED">
      <CLUB name="Feijenoord Albion Zwemclub" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:33.26">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-02" nation="NED" />
     <RELAY name="ZPC DE HOF" nation="NED">
      <CLUB name="ZPC DE HOF" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jasper" nameprefix="de" lastname="Boer" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Pieter" nameprefix="" lastname="Pickhardt" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Emiel" nameprefix="" lastname="Huisken" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Huisken" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:34.34">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Gwangju" date="2019-08-16" nation="KOR" />
     <RELAY name="Getxo" nation="ESP">
      <CLUB name="Getxo" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:43.83">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Kazan" date="2015-08-14" nation="RUS" />
     <RELAY name="Troyka Moscow" nation="RUS">
      <CLUB name="Troyka Moscow" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:33.25">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Riccione" date="2019-12-07" nation="ITA" />
     <RELAY name="Maranello Nuoto" nation="ITA">
      <CLUB name="Maranello Nuoto" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:58.35">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Kazan" date="2015-04-17" nation="RUS" />
     <RELAY name="Troyka Moscow" nation="RUS">
      <CLUB name="Troyka Moscow" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:56.92">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="St. Petersburg" date="2022-07-27" nation="RUS" />
     <RELAY name="Tsunami Nizhniy" nation="RUS">
      <CLUB name="Tsunami Nizhniy" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:31.95">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2009-11-29" nation="" />
     <RELAY name="MAC-MINA" nation="BRA">
      <CLUB name="MAC-MINA" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rene" nameprefix="" lastname="Leite" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rodrigo" nameprefix="" lastname="Trivino" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Daniel" nameprefix="" lastname="Belini" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Piero" nameprefix="" lastname="Rodigheri" gender="M" nation="BRA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:41.78">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-09-03" nation="" />
     <RELAY name="JFE Keihin" nation="JPN">
      <CLUB name="JFE Keihin" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:30.77">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2013-06-23" nation="" />
     <RELAY name="G-TRAVELERS" nation="JPN">
      <CLUB name="G-TRAVELERS" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Yoshinori" nameprefix="" lastname="Muramatsu" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kosuke" nameprefix="" lastname="Maeda" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Kensuke" nameprefix="" lastname="Maeda" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Naofumi" nameprefix="" lastname="Utsugi" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:46.80">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-09-19" nation="" />
     <RELAY name="Mitsuuroko" nation="JPN">
      <CLUB name="Mitsuuroko" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:39.05">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-09-03" nation="" />
     <RELAY name="JFE Keihin" nation="JPN">
      <CLUB name="JFE Keihin" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:40.52">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Londen" date="2016-05-26" nation="GBR" />
     <RELAY name="d&apos;ELFT" nation="NED">
      <CLUB name="d&apos;ELFT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Roderik" nameprefix="" lastname="Meijers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:51.61">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Londen" date="2016-05-27" nation="GBR" />
     <RELAY name="d&apos;ELFT WAVE (SG)" nation="NED">
      <CLUB name="d&apos;ELFT WAVE (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Egbert" nameprefix="" lastname="Stolk" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Simons" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Roderik" nameprefix="" lastname="Meijers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:45.50">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <RELAY name="Blue Marlins" nation="NED">
      <CLUB name="Blue Marlins" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jonne" nameprefix="" lastname="Schaafsma" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Stefan" nameprefix="" lastname="Petersen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jim" nameprefix="" lastname="Geestman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:04.86">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2017-05-07" nation="NED" />
     <RELAY name="Albion d&apos;ELFT (SG)" nation="NED">
      <CLUB name="Albion d&apos;ELFT (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ensger" nameprefix="" lastname="Kotterink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Romero" nameprefix="" lastname="Hennep" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Hugo" nameprefix="" lastname="Bregman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:39.33">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-02" nation="NED" />
     <RELAY name="Zwemlust-den Hommel" nation="NED">
      <CLUB name="Zwemlust-den Hommel" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Vincent" nameprefix="" lastname="Versteeg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Mark" nameprefix="" lastname="Musch" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Mark" nameprefix="" lastname="Zwart" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Raoul" nameprefix="" lastname="Engelenburg" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:32.84">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Reus" date="2018-07-08" nation="ESP" />
     <RELAY name="GETXO" nation="ESP">
      <CLUB name="GETXO" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:43.35">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2021-04-17" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novgorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novgorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:28.93">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Reus" date="2018-07-07" nation="ESP" />
     <RELAY name="GETXO" nation="ESP">
      <CLUB name="GETXO" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:58.88">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Serravalle" date="2023-05-06" nation="SMA" />
     <RELAY name="Amici Nuoto Firenze" nation="ITA">
      <CLUB name="Amici Nuoto Firenze" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:02.91">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Serravalle" date="2023-05-06" nation="SMA" />
     <RELAY name="Amici Nuoto Firenze" nation="ITA">
      <CLUB name="Amici Nuoto Firenze" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:32.84">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2018-07-08" nation="" />
     <RELAY name="GETXO" nation="ESP">
      <CLUB name="GETXO" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Mikel" nameprefix="" lastname="Bildosola Agirregomezkorta" gender="M" nation="ESP" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Inaki" nameprefix="" lastname="Bildosola" gender="M" nation="ESP" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="German" nameprefix="" lastname="Zubiaur" gender="M" nation="ESP" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Mikel" nameprefix="" lastname="Deba" gender="M" nation="ESP" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:42.06">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-05-27" nation="" />
     <RELAY name="CSKA" nation="RUS">
      <CLUB name="CSKA" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:28.93">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2018-07-07" nation="" />
     <RELAY name="GETXO" nation="ESP">
      <CLUB name="GETXO" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Mikel" nameprefix="" lastname="Bildosola Agirregomezkorta" gender="M" nation="ESP" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Inaki" nameprefix="" lastname="Bildosola" gender="M" nation="ESP" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="German" nameprefix="" lastname="Zubiaur" gender="M" nation="ESP" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Mikel" nameprefix="" lastname="Deba" gender="M" nation="ESP" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:49.75">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2019-01-19" nation="" />
     <RELAY name="JFE KEIHIN" nation="JPN">
      <CLUB name="JFE KEIHIN" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Takashi" nameprefix="" lastname="Takemoto" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hajime" nameprefix="" lastname="Ikegami" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ryoya" nameprefix="" lastname="Taguchi" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Shintaro" nameprefix="" lastname="Uchiyama" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:50.34">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-08-19" nation="" />
     <RELAY name="JFE" nation="JPN">
      <CLUB name="JFE" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ryoya" nameprefix="" lastname="Taguchi" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Takashi" nameprefix="" lastname="Takemoto" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Shintaro" nameprefix="" lastname="Uchiyama" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Takao" nameprefix="" lastname="Ueki" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:43.25">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Dennis" nameprefix="" lastname="Bos" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ren�" nameprefix="" lastname="Beetsma" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:56.93">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ren�" nameprefix="" lastname="Beetsma" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Dennis" nameprefix="" lastname="Bos" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:51.14">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Dennis" nameprefix="" lastname="Bos" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ren�" nameprefix="" lastname="Beetsma" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:18.44">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Alkmaar" date="2019-04-14" nation="NED" />
     <RELAY name="DAW" nation="NED">
      <CLUB name="DAW" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jorrick" nameprefix="" lastname="Druyven" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Joost" nameprefix="" lastname="Hoetjes" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Pieter" nameprefix="van" lastname="Gemeren" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Alex" nameprefix="" lastname="Damen" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:47.18">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Dennis" nameprefix="" lastname="Bos" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ren�" nameprefix="" lastname="Beetsma" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:34.92">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Neva Stars St Petersburg" nation="RUS">
      <CLUB name="Neva Stars St Petersburg" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Aleksandr" nameprefix="" lastname="Shilin" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:45.47">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Neva Stars St Petersburg" nation="RUS">
      <CLUB name="Neva Stars St Petersburg" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:39.87">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Brescia" date="2018-05-13" nation="ITA" />
     <RELAY name="AICS Aquare Mafeco" nation="ITA">
      <CLUB name="AICS Aquare Mafeco" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:02.57">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Brescia" date="2015-05-17" nation="ITA" />
     <RELAY name="Master AICS Brescia" nation="ITA">
      <CLUB name="Master AICS Brescia" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:11.34">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Brescia" date="2015-05-15" nation="ITA" />
     <RELAY name="Master AICS Bescia" nation="ITA">
      <CLUB name="Master AICS Bescia" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:34.92">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-08-18" nation="" />
     <RELAY name="NEVA STARS" nation="RUS">
      <CLUB name="NEVA STARS" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Aleksandr" nameprefix="" lastname="Shilin" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Sergei" nameprefix="" lastname="Medvedev" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Aleksei" nameprefix="" lastname="Manzhula" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Vladimir" nameprefix="" lastname="Predkin" gender="M" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:45.47">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-08-18" nation="" />
     <RELAY name="NEVA STARS" nation="RUS">
      <CLUB name="NEVA STARS" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Aleksandr" nameprefix="" lastname="Shilin" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Sergey" nameprefix="" lastname="Gogol" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Aleksei" nameprefix="" lastname="Manzhula" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Vladimir" nameprefix="" lastname="Predkin" gender="M" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:38.60">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2011-07-03" nation="" />
     <RELAY name="LONGHORN AQUATICS" nation="USA">
      <CLUB name="LONGHORN AQUATICS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Tyler" nameprefix="" lastname="Blessing" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Mike" nameprefix="" lastname="Varozza" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anders" nameprefix="" lastname="Rasmussen" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Chris" nameprefix="" lastname="Eckerman" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:01.27">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-03-12" nation="" />
     <RELAY name="Diablo" nation="JPN">
      <CLUB name="Diablo" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:12.71">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-10-24" nation="" />
     <RELAY name="JSS Fukai" nation="JPN">
      <CLUB name="JSS Fukai" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:48.09">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <RELAY name="AZ&amp;PC De Futen" nation="NED">
      <CLUB name="AZ&amp;PC De Futen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Gert" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Bas" nameprefix="" lastname="Tappel" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Arnold" nameprefix="de" lastname="Rover" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Dennis" nameprefix="" lastname="Kos" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:00.63">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jeroen" nameprefix="" lastname="Zelsmann" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:03.54">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-06" nation="NED" />
     <RELAY name="De Rog" nation="NED">
      <CLUB name="De Rog" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Arjan" nameprefix="" lastname="Verheij" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Spetter" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Glen" nameprefix="le" lastname="Clercq" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:48.44">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <RELAY name="De Rog" nation="NED">
      <CLUB name="De Rog" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Kamphuis" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Glen" nameprefix="le" lastname="Clercq" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Spetter" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:26.96">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2016-05-06" nation="NED" />
     <RELAY name="De Rog" nation="NED">
      <CLUB name="De Rog" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Spetter" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Kamphuis" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Glen" nameprefix="le" lastname="Clercq" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:41.19">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Riccione" date="2016-06-26" nation="ITA" />
     <RELAY name="Centro Nuoto Bastilia" nation="ITA">
      <CLUB name="Centro Nuoto Bastilia" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:52.36">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Nuoto Masters Brescia" nation="ITA">
      <CLUB name="Nuoto Masters Brescia" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:46.05">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Lamarmora" date="2017-05-14" nation="ITA" />
     <RELAY name="AICS Acquare Mafeco" nation="ITA">
      <CLUB name="AICS Acquare Mafeco" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:14.38">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Brescia" date="2017-05-13" nation="ITA" />
     <RELAY name="Brescia Acquare Mafeco" nation="ITA">
      <CLUB name="Brescia Acquare Mafeco" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:47.63">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <RELAY name="Oslo Idrettslag Sv�mming" nation="NOR">
      <CLUB name="Oslo Idrettslag Sv�mming" nation="NOR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="�ivind Martin" nameprefix="" lastname="Hasle" gender="M" nation="NOR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Knut Ivan" nameprefix="" lastname="Rasmussen" gender="M" nation="NOR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erlend" nameprefix="" lastname="Alstad" gender="M" nation="NOR" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Oddvar" nameprefix="" lastname="Sandvin" gender="M" nation="NOR" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:38.24">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2006-08-08" nation="" />
     <RELAY name="COLORADO MASTERS" nation="USA">
      <CLUB name="COLORADO MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jack" nameprefix="" lastname="Groselle" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Trip" nameprefix="" lastname="Hedrick" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Steve" nameprefix="" lastname="Wood" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:50.83">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2006-08-08" nation="" />
     <RELAY name="COLORADO MASTERS" nation="USA">
      <CLUB name="COLORADO MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Steve" nameprefix="" lastname="Wood" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jack" nameprefix="" lastname="Groselle" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Trip" nameprefix="" lastname="Hedrick" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:46.05">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-05-14" nation="" />
     <RELAY name="BRESCIA ACQUARE MAFECO" nation="ITA">
      <CLUB name="BRESCIA ACQUARE MAFECO" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Massimiliano" nameprefix="" lastname="Gialdi" gender="M" nation="ITA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Maurizio" nameprefix="" lastname="Tersar" gender="M" nation="ITA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Roberto" nameprefix="" lastname="Brunori" gender="M" nation="ITA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marco" nameprefix="" lastname="Colombo" gender="M" nation="ITA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:13.76">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2012-08-11" nation="" />
     <RELAY name="LONGHORN AQUATICS" nation="USA">
      <CLUB name="LONGHORN AQUATICS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Anders" nameprefix="" lastname="Rasmussen" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jim" nameprefix="" lastname="Sauer" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="David" nameprefix="" lastname="Guthrie" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Mike" nameprefix="" lastname="Varozza" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:38.24">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2013-07-06" nation="" />
     <RELAY name="BRASIL MASTERS" nation="BRA">
      <CLUB name="BRASIL MASTERS" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Helio" nameprefix="" lastname="Celidonio" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Djan" nameprefix="" lastname="Garrido Madruga" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Roberto Carlos" nameprefix="" lastname="Carvalho" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marcus" nameprefix="" lastname="Mattioli" gender="M" nation="BRA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:54.53">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-07" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Joop" nameprefix="" lastname="Ariaens" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:11.97">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2017-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Joop" nameprefix="" lastname="Ariaens" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:17.68">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Joop" nameprefix="" lastname="Ariaens" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:56.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Harold" nameprefix="" lastname="Matla" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:20.84">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <RELAY name="De Rog" nation="NED">
      <CLUB name="De Rog" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Kamphuis" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Roy" nameprefix="le" lastname="Clercq" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Spetter" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Peter" nameprefix="" lastname="Bernsen" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:49.16">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Goeteborg" nation="SWE">
      <CLUB name="Goeteborg" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Leonard" nameprefix="" lastname="Bielicz" gender="M" nation="SWE" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:03.70">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="G�teborg Sim" nation="DEN">
      <CLUB name="G�teborg Sim" nation="DEN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:17.68">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Joop" nameprefix="" lastname="Ariaens" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:51.54">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Las Palmas" date="2023-06-19" nation="ESP" />
     <RELAY name="Tenerife Masters" nation="ESP">
      <CLUB name="Tenerife Masters" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:42.09">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="St. Petersburg" date="2022-04-24" nation="RUS" />
     <RELAY name="Tsunami Nizhniy" nation="RUS">
      <CLUB name="Tsunami Nizhniy" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:42.40">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2016-08-19" nation="" />
     <RELAY name="SARASOTA Y SHARKS" nation="USA">
      <CLUB name="SARASOTA Y SHARKS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Steve" nameprefix="" lastname="Wood" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Doug" nameprefix="" lastname="Martin" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Trip" nameprefix="" lastname="Hedrick" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jack" nameprefix="" lastname="Groselle" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:57.46">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-08-21" nation="" />
     <RELAY name="SARASOTA Y SHARKS" nation="USA">
      <CLUB name="SARASOTA Y SHARKS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Steve" nameprefix="" lastname="Wood" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jack" nameprefix="" lastname="Groselle" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Trip" nameprefix="" lastname="Hedrick" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Doug" nameprefix="" lastname="Martin" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:59.86">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2018-08-11" nation="" />
     <RELAY name="COLORADO MASTERS" nation="USA">
      <CLUB name="COLORADO MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Craig" nameprefix="" lastname="Petersen" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Greg" nameprefix="" lastname="Scott" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Kirk" nameprefix="" lastname="Anderson" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:32.15">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2018-08-10" nation="" />
     <RELAY name="COLORADO MASTERS" nation="USA">
      <CLUB name="COLORADO MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Craig" nameprefix="" lastname="Petersen" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Greg" nameprefix="" lastname="Scott" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Kirk" nameprefix="" lastname="Anderson" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:56.62">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2018-08-12" nation="" />
     <RELAY name="COLORADO MASTERS" nation="USA">
      <CLUB name="COLORADO MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Michael" nameprefix="" lastname="Mann" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Craig" nameprefix="" lastname="Petersen" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Greg" nameprefix="" lastname="Scott" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Kirk" nameprefix="" lastname="Anderson" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:21.93">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jan" nameprefix="" lastname="Tinholt" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:47.15">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hemesath" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jan" nameprefix="" lastname="Nuijten" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:39.85">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Fred" nameprefix="" lastname="Ketting" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jan" nameprefix="" lastname="Nuijten" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Andr�" nameprefix="" lastname="Pantekoek" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:17.00">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Ron" nameprefix="" lastname="Phaff" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:12:44.37">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Hans" nameprefix="" lastname="Wijsman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:00.76">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Vichy" date="2009-06-13" nation="FRA" />
     <RELAY name="CN MARSEILLE" nation="FRA">
      <CLUB name="CN MARSEILLE" nation="FRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:18.10">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Totokbalinti Senior" nation="HUN">
      <CLUB name="Totokbalinti Senior" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:46.27">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Ravenna" date="2020-01-12" nation="ITA" />
     <RELAY name="DLF Nuoto Livorno" nation="ITA">
      <CLUB name="DLF Nuoto Livorno" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:37.43">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2012-05-05" nation="GBR" />
     <RELAY name="BIRMINGHAM MASTERS" nation="GBR">
      <CLUB name="BIRMINGHAM MASTERS" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:11:07.44">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Las Palmas" date="2023-06-19" nation="ESP" />
     <RELAY name="Tenerife Masters" nation="ESP">
      <CLUB name="Tenerife Masters" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:53.43">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-08-05" nation="" />
     <RELAY name="Swim Fort Lauderdale" nation="USA">
      <CLUB name="Swim Fort Lauderdale" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:07.03">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-08-04" nation="" />
     <RELAY name="Swim Fort Lauderdale" nation="USA">
      <CLUB name="Swim Fort Lauderdale" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:27.17">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-06-18" nation="" />
     <RELAY name="PALM BEACH MASTERS" nation="USA">
      <CLUB name="PALM BEACH MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lee" nameprefix="" lastname="Childs" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Keefe" nameprefix="" lastname="Lodwig" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="George" nameprefix="" lastname="Schmidt" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="David" nameprefix="" lastname="Quiggin" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:07.90">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-08-07" nation="" />
     <RELAY name="Saratosa Sharks" nation="USA">
      <CLUB name="Saratosa Sharks" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:15.72">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-06-06" nation="" />
     <RELAY name="SARASOTA SHARKS" nation="USA">
      <CLUB name="SARASOTA SHARKS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jack" nameprefix="" lastname="Groselle" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Couch" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Rick" nameprefix="" lastname="Walker" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:26.67">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Kranj" date="2018-09-05" nation="SLO" />
     <RELAY name="Hellas" nation="SWE">
      <CLUB name="Hellas" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Erik" nameprefix="" lastname="Forslund" gender="M" nation="SWE" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Anders" nameprefix="" lastname="S�derqvist" gender="M" nation="SWE" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Peter" nameprefix="" lastname="Bergengren" gender="M" nation="SWE" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:48.59">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Gyula" date="2023-06-23" nation="HUN" />
     <RELAY name="T�r�kb�lint Senior" nation="HUN">
      <CLUB name="T�r�kb�lint Senior" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:09.75">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Magdeburg" date="2017-06-16" nation="GER" />
     <RELAY name="SSV Leutsch Leipzig" nation="GER">
      <CLUB name="SSV Leutsch Leipzig" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:40.23">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Kecskemet" date="2023-04-15" nation="HUN" />
     <RELAY name="T�r�kb�lint Senior" nation="HUN">
      <CLUB name="T�r�kb�lint Senior" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:13:47.68">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Dresden" date="2017-05-06" nation="GER" />
     <RELAY name="SSV Leutsch Leipzig" nation="GER">
      <CLUB name="SSV Leutsch Leipzig" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:12.73">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-07-23" nation="" />
     <RELAY name="Tamalpais Aquatic Masters" nation="USA">
      <CLUB name="Tamalpais Aquatic Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:37.00">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-07-22" nation="" />
     <RELAY name="Tamalpais Aquatic Masters" nation="USA">
      <CLUB name="Tamalpais Aquatic Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:05.88">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-07-22" nation="" />
     <RELAY name="Tamalpais Aquatic Masters" nation="USA">
      <CLUB name="Tamalpais Aquatic Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:14.23">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-07-23" nation="" />
     <RELAY name="Tamalpais Aquatic  Masters" nation="USA">
      <CLUB name="Tamalpais Aquatic  Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:11:38.85">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-07-21" nation="" />
     <RELAY name="Tamalpais Aquatic Masters" nation="USA">
      <CLUB name="Tamalpais Aquatic Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:04:57.70">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Gavrylych Swim Club" nation="UKR">
      <CLUB name="Gavrylych Swim Club" nation="UKR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:26.29">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Gavrylych Swim Club" nation="UKR">
      <CLUB name="Gavrylych Swim Club" nation="UKR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:56.10">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Zaporizhzhiya" date="2017-03-25" nation="UKR" />
     <RELAY name="Gavrylych SC" nation="UKR">
      <CLUB name="Gavrylych SC" nation="UKR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:12:23.62">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Dnipro" date="2017-05-13" nation="UKR" />
     <RELAY name="Gavryilych swim club" nation="UKR">
      <CLUB name="Gavryilych swim club" nation="UKR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="M" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:03:08.87">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2008-03-02" nation="" />
     <RELAY name="JUEI CLUB" nation="JPN">
      <CLUB name="JUEI CLUB" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Isamu" nameprefix="" lastname="Tamura" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Tokushi" nameprefix="" lastname="Komeda" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Hideya" nameprefix="" lastname="Fujii" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Hidekazu" nameprefix="" lastname="Tamura" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:13.40">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2009-06-20" nation="" />
     <RELAY name="NISHINOMIYA SUMIRE" nation="JPN">
      <CLUB name="NISHINOMIYA SUMIRE" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Roshio" nameprefix="" lastname="Yuri" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Takeshi" nameprefix="" lastname="Yasukawa" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Himoru" nameprefix="" lastname="Yoshimoto" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Kazunaga" nameprefix="" lastname="Akutsu" gender="M" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:03.44">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-07-10" nation="" />
     <RELAY name="San Diego Masters swimming" nation="USA">
      <CLUB name="San Diego Masters swimming" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:11:32.00">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-04-30" nation="" />
     <RELAY name="Victor Spiritus Power" nation="BRA">
      <CLUB name="Victor Spiritus Power" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:24:45.07">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-04-30" nation="" />
     <RELAY name="Victor Spiritus Power" nation="BRA">
      <CLUB name="Victor Spiritus Power" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="80" agemax="99" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:44.27">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-04" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Kimberley" nameprefix="" lastname="Albers" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Anja" nameprefix="van der" lastname="Hout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Bruno" nameprefix="" lastname="Carissimi Boff" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Mark" nameprefix="" lastname="Costeris" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:57.14">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2014-05-03" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Anja" nameprefix="van der" lastname="Hout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Isabelle" nameprefix="" lastname="Massar" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Bruno" nameprefix="" lastname="Carissimi Boff" gender="M" nation="BRA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Mark" nameprefix="" lastname="Costeris" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:55.20">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="Nova" nation="NED">
      <CLUB name="Nova" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Roy" nameprefix="" lastname="Smeenge" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lisanne" nameprefix="" lastname="Boets" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Karin" nameprefix="" lastname="Groen" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Darren" nameprefix="" lastname="Chen" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:22.90">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <RELAY name="ZVL-1886 Center" nation="NED">
      <CLUB name="ZVL-1886 Center" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Sanne" nameprefix="" lastname="Heemskerk" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Silke" nameprefix="" lastname="Molendijk" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Robin" nameprefix="van" lastname="Beek" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Guus" nameprefix="" lastname="Hoogduin" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:50.88">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <RELAY name="ZVL-1886 Center" nation="NED">
      <CLUB name="ZVL-1886 Center" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Guus" nameprefix="" lastname="Hoogduin" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Robin" nameprefix="van" lastname="Beek" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Karen" nameprefix="" lastname="Stolk" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Silke" nameprefix="" lastname="Molendijk" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:41.21">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-09-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rieneke" nameprefix="" lastname="Terink" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Geert" nameprefix="" lastname="Lantink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjolijn" nameprefix="" lastname="Wuisman" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Stefan" nameprefix="" lastname="Oosting" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:53.92">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="Blue Marlins (SG)" nation="NED">
      <CLUB name="Blue Marlins (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Babette" nameprefix="van der" lastname="Kaaij" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Stefan" nameprefix="" lastname="Petersen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ilse" nameprefix="" lastname="Kraaijeveld" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:55.04">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="Blue Marlins (SG)" nation="NED">
      <CLUB name="Blue Marlins (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jim" nameprefix="" lastname="Geestman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Myra" nameprefix="" lastname="Smulders" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jeroen" nameprefix="" lastname="Baars" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Ilse" nameprefix="" lastname="Kraaijeveld" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:22.53">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2013-05-04" nation="NED" />
     <RELAY name="ZWEMLUST-DEN HOMMEL" nation="NED">
      <CLUB name="ZWEMLUST-DEN HOMMEL" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Charlotte" nameprefix="" lastname="Groeneveld" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Vincent" nameprefix="" lastname="Versteeg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Sven" nameprefix="" lastname="Jaeger" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Malissa" nameprefix="van der" lastname="Horst" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:44.61">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2017-05-05" nation="NED" />
     <RELAY name="WVZ" nation="NED">
      <CLUB name="WVZ" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Delia" nameprefix="" lastname="Badoux" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Isabelle" nameprefix="" lastname="Massar" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Bryan" nameprefix="" lastname="Mannaart" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Rutger" nameprefix="van" lastname="Oosterhout" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:41.21">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2013-09-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rieneke" nameprefix="" lastname="Terink" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Geert" nameprefix="" lastname="Lantink" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjolijn" nameprefix="" lastname="Wuisman" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Stefan" nameprefix="" lastname="Oosting" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:52.57">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Kazan" date="2015-08-14" nation="RUS" />
     <RELAY name="Poseidon Moscow" nation="RUS">
      <CLUB name="Poseidon Moscow" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:48.68">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Hannover" date="2014-06-20" nation="GER" />
     <RELAY name="W98 HANNOVER" nation="GER">
      <CLUB name="W98 HANNOVER" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Tim" nameprefix="" lastname="Grabowski" gender="M" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Constantin" nameprefix="" lastname="Dahle" gender="M" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anna Sophie" nameprefix="" lastname="Marx" gender="F" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nina-Christin" nameprefix="" lastname="Winter" gender="F" nation="GER" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:16.68">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:39.12">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Vitoria" date="2019-04-27" nation="ESP" />
     <RELAY name="Monteverde" nation="ESP">
      <CLUB name="Monteverde" nation="ESP" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="100" agemax="119" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:38.55">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-06-24" nation="" />
     <RELAY name="Swim Easy SPB" nation="RUS">
      <CLUB name="Swim Easy SPB" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:47.29">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-06-25" nation="" />
     <RELAY name="Swim-Easy SPB" nation="RUS">
      <CLUB name="Swim-Easy SPB" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:48.68">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Hannover" date="2014-06-20" nation="GER" />
     <RELAY name="W98 HANNOVER" nation="GER">
      <CLUB name="W98 HANNOVER" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Tim" nameprefix="" lastname="Grabowski" gender="M" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Constantin" nameprefix="" lastname="Dahle" gender="M" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Anna Sophie" nameprefix="" lastname="Marx" gender="F" nation="GER" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nina-Christin" nameprefix="" lastname="Winter" gender="F" nation="GER" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:05.01">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-03-12" nation="" />
     <RELAY name="Queendom" nation="JPN">
      <CLUB name="Queendom" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:35.56">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2019-12-15" nation="" />
     <RELAY name="SEN-SWIM" nation="JPN">
      <CLUB name="SEN-SWIM" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Tomoki" nameprefix="" lastname="Tanaka" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Chikahide" nameprefix="" lastname="Endo" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Kanako" nameprefix="" lastname="Tayama" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Mikiko" nameprefix="" lastname="Ito" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:42.44">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2004-02-15" nation="NED" />
     <RELAY name="AZ&amp;PC" nation="NED">
      <CLUB name="AZ&amp;PC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Annabel" nameprefix="" lastname="Kosten" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Tamara" nameprefix="van" lastname="Gorkom" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:57.54">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Martijn" nameprefix="" lastname="Giezen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:00.28">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-08" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jan-Willem" nameprefix="van der" lastname="Graaff" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Soraya" nameprefix="" lastname="Wasser" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Nelly" nameprefix="" lastname="Velthuijs" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Youri" nameprefix="" lastname="Vaes" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:23.51">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Martijn" nameprefix="" lastname="Giezen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:53.72">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <RELAY name="Albion d&apos;ELFT (SG)" nation="NED">
      <CLUB name="Albion d&apos;ELFT (SG)" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Timo" nameprefix="" lastname="Dinkelberg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Roos" nameprefix="van" lastname="Esch" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Dinkelberg" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nol" nameprefix="van" lastname="Thull" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:40.14">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Kazan" date="2015-08-14" nation="RUS" />
     <RELAY name="Tsunami Nizhniy Novgorod" nation="RUS">
      <CLUB name="Tsunami Nizhniy Novgorod" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:51.75">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Saransk" date="2021-04-18" nation="RUS" />
     <RELAY name="Tsunami" nation="RUS">
      <CLUB name="Tsunami" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:52.56">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Saransk" date="2021-04-17" nation="RUS" />
     <RELAY name="Lada Tolvatti" nation="RUS">
      <CLUB name="Lada Tolvatti" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:15.05">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Serravalle" date="2022-05-08" nation="ITA" />
     <RELAY name="Roma Nuoto Masters" nation="ITA">
      <CLUB name="Roma Nuoto Masters" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:25.05">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-02" nation="GBR" />
     <RELAY name="Trafford Metro" nation="GBR">
      <CLUB name="Trafford Metro" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="120" agemax="159" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:40.14">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-08-14" nation="" />
     <RELAY name="TSUNAMI" nation="RUS">
      <CLUB name="TSUNAMI" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Alexandr" nameprefix="" lastname="Satanovskiy" gender="M" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Irina" nameprefix="" lastname="Shlemova" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Svetlana" nameprefix="" lastname="Kniaginina" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Andrey" nameprefix="" lastname="Krylov" gender="M" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:49.61">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-05-28" nation="" />
     <RELAY name="Tusnami" nation="RUS">
      <CLUB name="Tusnami" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:49.88">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-10-07" nation="" />
     <RELAY name="Portiguar Masters" nation="BRA">
      <CLUB name="Portiguar Masters" nation="BRA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:14.85">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-09-17" nation="" />
     <RELAY name="Frontier RC" nation="JPN">
      <CLUB name="Frontier RC" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:25.05">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-06-02" nation="" />
     <RELAY name="Trafford Met" nation="GBR">
      <CLUB name="Trafford Met" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:48.90">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Millau" date="2003-08-29" nation="FRA" />
     <RELAY name="AZ&amp;PC" nation="NED">
      <CLUB name="AZ&amp;PC" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Petra" nameprefix="" lastname="Casteleijn-Frowijn" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Peter" nameprefix="van" lastname="Meerveld" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:00.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Martijn" nameprefix="" lastname="Giezen" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Larissa" nameprefix="" lastname="Brak" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:06.63">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Danielle" nameprefix="de" lastname="Boer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:38.28">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2022-05-07" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jelle" nameprefix="" lastname="Opmeer" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marije" nameprefix="" lastname="Jansen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:18.16">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-01-06" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ren�" nameprefix="" lastname="Beetsma" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Danielle" nameprefix="de" lastname="Boer" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Casper" nameprefix="" lastname="Hut" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:42.77">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="St. Petersburg" date="2015-06-07" nation="RUS" />
     <RELAY name="Neva Stars St.Petersburg" nation="RUS">
      <CLUB name="Neva Stars St.Petersburg" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:55.32">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Kazan" date="2015-08-14" nation="RUS" />
     <RELAY name="Neva Stars-St.Petersburg" nation="RUS">
      <CLUB name="Neva Stars-St.Petersburg" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:56.44">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Szentes" date="2017-01-21" nation="HUN" />
     <RELAY name="Iron Aquatics" nation="HUN">
      <CLUB name="Iron Aquatics" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:21.61">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Swansea" date="2019-06-14" nation="GBR" />
     <RELAY name="Fareham Nomads" nation="GBR">
      <CLUB name="Fareham Nomads" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:44.02">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Brescia" date="2019-05-12" nation="ITA" />
     <RELAY name="Nuoto Master Brescia" nation="ITA">
      <CLUB name="Nuoto Master Brescia" nation="ITA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="160" agemax="199" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:42.27">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2006-08-08" nation="" />
     <RELAY name="TEAM TYR" nation="USA">
      <CLUB name="TEAM TYR" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="John" nameprefix="" lastname="Smith" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Saeger" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Collette" nameprefix="" lastname="Sappey" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Sheri" nameprefix="" lastname="Hart" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:53.25">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2021-06-06" nation="" />
     <RELAY name="Mad Wave" nation="RUS">
      <CLUB name="Mad Wave" nation="RUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Alexandra" nameprefix="" lastname="Povaliy" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Anna" nameprefix="" lastname="Polyakova" gender="F" nation="RUS" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Vladislav" nameprefix="" lastname="Bragin" gender="M" nation="CZE" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Vladimir" nameprefix="" lastname="Predkin" gender="M" nation="RUS" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:51.77">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-12-02" nation="" />
     <RELAY name="CBH" nation="PAR">
      <CLUB name="CBH" nation="PAR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:15.64">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-06-18" nation="" />
     <RELAY name="JSS Fukai" nation="JPN">
      <CLUB name="JSS Fukai" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:43.94">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-11-11" nation="" />
     <RELAY name="BP HONVED SE" nation="HUN">
      <CLUB name="BP HONVED SE" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Melinda" nameprefix="" lastname="Marosi" gender="F" nation="HUN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Dora" nameprefix="" lastname="Cerva" gender="F" nation="HUN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Andras" nameprefix="" lastname="Schonek" gender="M" nation="HUN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Valter" nameprefix="" lastname="Kalaus" gender="M" nation="HUN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:51.50">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Jeroen" nameprefix="" lastname="Zelsmann" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:07.81">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Vincent" nameprefix="" lastname="Bakker" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:15.97">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-04" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Erwin" nameprefix="" lastname="Buist" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:46.35">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2019-05-05" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Vincent" nameprefix="" lastname="Bakker" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lesley" nameprefix="" lastname="Cordial" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:46.40">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2019-05-03" nation="NED" />
     <RELAY name="HZ&amp;PC Heerenveen" nation="NED">
      <CLUB name="HZ&amp;PC Heerenveen" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Ren�" nameprefix="" lastname="Beetsma" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jannie" nameprefix="" lastname="Vennik" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Evelien" nameprefix="van" lastname="Klaarbergen-Kleinhuis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Marten" nameprefix="de" lastname="Groot" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:47.37">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Berliner TSC" nation="GER">
      <CLUB name="Berliner TSC" nation="GER" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Budapest" date="2017-08-18" nation="HUN" />
     <RELAY name="Guildford City Swim" nation="GBR">
      <CLUB name="Guildford City Swim" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:05.39">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <RELAY name="Woking" nation="GBR">
      <CLUB name="Woking" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:33.51">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Sheffield" date="2023-06-03" nation="GBR" />
     <RELAY name="Woking" nation="GBR">
      <CLUB name="Woking" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:12.43">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Sheffield" date="2023-06-02" nation="GBR" />
     <RELAY name="Woking" nation="GBR">
      <CLUB name="Woking" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="200" agemax="239" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:44.96">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2006-08-08" nation="" />
     <RELAY name="COLORADO MASTERS" nation="USA">
      <CLUB name="COLORADO MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Trip" nameprefix="" lastname="Hedrick" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kim" nameprefix="" lastname="Crouch" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Kathy" nameprefix="" lastname="Garnier" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Abrahams" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:01:57.86">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-08-05" nation="" />
     <RELAY name="North Carolina Masters" nation="USA">
      <CLUB name="North Carolina Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:57.74">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-05-07" nation="" />
     <RELAY name="Powerpoints" nation="AUS">
      <CLUB name="Powerpoints" nation="AUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:30.56">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2023-08-20" nation="" />
     <RELAY name="North Carolina Masters" nation="USA">
      <CLUB name="North Carolina Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:55.03">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-03-03" nation="" />
     <RELAY name="Powerpoints" nation="AUS">
      <CLUB name="Powerpoints" nation="AUS" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:56.14">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:08.71">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:20.39">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:00.59">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:44.46">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:56.14">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:08.71">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:20.39">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-06" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Edwin" nameprefix="van" lastname="Norden" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:52.45">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Aberdeen" date="2022-06-17" nation="GBR" />
     <RELAY name="Spencer" nation="GBR">
      <CLUB name="Spencer" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:44.46">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Amersfoort" date="2023-05-05" nation="NED" />
     <RELAY name="ZPC AMERSFOORT" nation="NED">
      <CLUB name="ZPC AMERSFOORT" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Chester" nameprefix="" lastname="Marsman" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Atie" nameprefix="" lastname="Pijtak-Radersma" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Marjan" nameprefix="" lastname="Remmits-de Lange" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Johan" nameprefix="" lastname="Remmits" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="240" agemax="279" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:01:54.54">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2016-08-20" nation="" />
     <RELAY name="SARASOTA Y SHARKS" nation="USA">
      <CLUB name="SARASOTA Y SHARKS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Doug" nameprefix="" lastname="Martin" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jack" nameprefix="" lastname="Groselle" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Nancy" nameprefix="" lastname="Kryka" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Laura" nameprefix="" lastname="Kirkpatrick" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:08.11">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2016-08-20" nation="" />
     <RELAY name="PUGET SOUND MASTERS" nation="USA">
      <CLUB name="PUGET SOUND MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lisa" nameprefix="" lastname="Dahl" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rick" nameprefix="" lastname="Colella" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Donald" nameprefix="" lastname="Graham" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Charlotte" nameprefix="" lastname="Davis" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:19.89">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2015-03-19" nation="" />
     <RELAY name="CAPE TOWN MASTERS" nation="RSA">
      <CLUB name="CAPE TOWN MASTERS" nation="RSA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Calvin" nameprefix="" lastname="Maughan" gender="M" nation="rsa" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Sanderina" nameprefix="" lastname="Kruger" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Diane" nameprefix="" lastname="Coetzee" gender="F" nation="RSA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Timothy" nameprefix="" lastname="Shead" gender="M" nation="RSA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:44.76">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2022-07-09" nation="" />
     <RELAY name="Lone star masters" nation="USA">
      <CLUB name="Lone star masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:35.54">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-07-22" nation="" />
     <RELAY name="Lone Star Masters" nation="USA">
      <CLUB name="Lone Star Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:23.07">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2014-05-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:45.76">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:11.01">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-05" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Brend" nameprefix="" lastname="Brev�" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Annie" nameprefix="" lastname="Smits" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Patty" nameprefix="" lastname="Verhagen" gender="F" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:35.90">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Amersfoort" date="2023-05-07" nation="NED" />
     <RELAY name="SWOL 1894" nation="NED">
      <CLUB name="SWOL 1894" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Berkhof" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Bea" nameprefix="" lastname="Swijnenberg" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Christine" nameprefix="" lastname="Nieuwenhuis" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Harry" nameprefix="" lastname="Dokter" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:13:57.75">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Den Haag" date="2018-05-04" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Katrin" nameprefix="" lastname="Pennings" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Annie" nameprefix="" lastname="Smits" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:14.78">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Fukuoka" date="2023-08-09" nation="JPN" />
     <RELAY name="Spencer Masters Swim Team" nation="GBR">
      <CLUB name="Spencer Masters Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:32.35">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Kranj" date="2018-09-04" nation="SLO" />
     <RELAY name="Torokbalitini Senior" nation="HUN">
      <CLUB name="Torokbalitini Senior" nation="HUN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Monika" nameprefix="" lastname="Balla" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="F" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="vacant" gender="M" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:20.02">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Crawley" date="2023-03-25" nation="GBR" />
     <RELAY name="Spencer Masters Swim Team" nation="GBR">
      <CLUB name="Spencer Masters Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:02.46">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Crawley" date="2023-03-25" nation="GBR" />
     <RELAY name="Spencer Masters Swim Team" nation="GBR">
      <CLUB name="Spencer Masters Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:11:39.59">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Crawley" date="2023-03-25" nation="GBR" />
     <RELAY name="Spencer Masters Swim Team" nation="GBR">
      <CLUB name="Spencer Masters Swim Team" nation="GBR" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="280" agemax="319" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:03.33">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2021-10-09" nation="" />
     <RELAY name="Tamalpais Aquatics" nation="USA">
      <CLUB name="Tamalpais Aquatics" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:21.20">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-08-09" nation="" />
     <RELAY name="TAMALPAIS AQUATIC MASTERS" nation="USA">
      <CLUB name="TAMALPAIS AQUATIC MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kenneth" nameprefix="" lastname="Frost" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nancy" nameprefix="" lastname="Ridout" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:45.34">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2023-07-09" nation="" />
     <RELAY name="Saratosa Sharks" nation="USA">
      <CLUB name="Saratosa Sharks" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:05:28.17">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2015-05-10" nation="" />
     <RELAY name="TAMALPAIS MASTERS" nation="USA">
      <CLUB name="TAMALPAIS MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Richard" nameprefix="" lastname="Burns" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Kenneth" nameprefix="" lastname="Frost" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Laura" nameprefix="" lastname="Val" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nancy" nameprefix="" lastname="Ridout" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:37.37">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-07-29" nation="" />
     <RELAY name="Tamalpais Masters" nation="USA">
      <CLUB name="Tamalpais Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:52.48">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Luxembourg/Hollerich" date="2021-10-10" nation="LUX" />
     <RELAY name="Psv" nation="NED">
      <CLUB name="Psv" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:34.35">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2017-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Wim" nameprefix="ter" lastname="Laak" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:16.29">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2015-05-09" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Cor" nameprefix="" lastname="Sprengers" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Bob" nameprefix="" lastname="Berg" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:09:21.81">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Eindhoven" date="2015-05-10" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Alice" nameprefix="" lastname="Lindhout" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Marianne" nameprefix="" lastname="Maandonks" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rob" nameprefix="" lastname="Hanou" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Cor" nameprefix="" lastname="Sprengers" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:15:16.47">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Eindhoven" date="2022-05-06" nation="NED" />
     <RELAY name="PSV" nation="NED">
      <CLUB name="PSV" nation="NED" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Corrie" nameprefix="" lastname="Verhoeven" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Lottie" nameprefix="" lastname="Geurts" gender="F" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jan" nameprefix="" lastname="Nuijten" gender="M" nation="NED" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Nic" nameprefix="" lastname="Geers" gender="M" nation="NED" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:52.02">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="Riccione" date="2004-06-08" nation="IRA" />
     <RELAY name="SOIK HELLAS" nation="SWE">
      <CLUB name="SOIK HELLAS" nation="SWE" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:03:04.72">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Charleroi" date="2016-04-17" nation="BEL" />
     <RELAY name="AZSC" nation="BEL">
      <CLUB name="AZSC" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:44.34">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="Wachtebeke" date="2016-02-27" nation="BEL" />
     <RELAY name="AZSC" nation="BEL">
      <CLUB name="AZSC" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:30.47">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="Charleroi" date="2016-04-17" nation="BEL" />
     <RELAY name="AZCS" nation="BEL">
      <CLUB name="AZCS" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:15:14.13">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="Charleroi" date="2016-04-16" nation="BEL" />
     <RELAY name="AZSC" nation="BEL">
      <CLUB name="AZSC" nation="BEL" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Agnes" nameprefix="" lastname="Van Obberghen-Pieters" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Eliane" nameprefix="" lastname="Pellis" gender="F" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jozef" nameprefix="van" lastname="Roy" gender="M" nation="BEL" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Joseph" nameprefix="" lastname="Meyten" gender="M" nation="BEL" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="320" agemax="359" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:02:35.97">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2016-08-20" nation="" />
     <RELAY name="OREGON MASTERS" nation="USA">
      <CLUB name="OREGON MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rebecca" nameprefix="" lastname="Kay" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Barbara" nameprefix="" lastname="Frid" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:02:55.98">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2014-07-20" nation="" />
     <RELAY name="BIG S YOKOHAMA" nation="JPN">
      <CLUB name="BIG S YOKOHAMA" nation="JPN" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Shoko" nameprefix="" lastname="Yonezawa" gender="F" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Hiyoshi" nameprefix="" lastname="Makimoto" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Tetsuo" nameprefix="" lastname="Nakamaru" gender="M" nation="JPN" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Meiko" nameprefix="" lastname="Kamashita" gender="F" nation="JPN" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:06:07.33">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2017-08-26" nation="" />
     <RELAY name="OREGON MASTERS" nation="USA">
      <CLUB name="OREGON MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Joy" nameprefix="" lastname="Ward" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Janet" nameprefix="" lastname="Gettling" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:07:17.49">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2017-08-27" nation="" />
     <RELAY name="OREGON MASTERS" nation="USA">
      <CLUB name="OREGON MASTERS" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Willard" nameprefix="" lastname="Lamb" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Ginger" nameprefix="" lastname="Pierson" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Joy" nameprefix="" lastname="Ward" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="David" nameprefix="" lastname="Radcliff" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:14:25.49">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2022-05-14" nation="" />
     <RELAY name="Oregon Masters" nation="USA">
      <CLUB name="Oregon Masters" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="NMR" name="Nederlands Masters Record" updated="2024-01-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="EMR" name="Europees Masters Record" updated="2023-11-30">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="23:59:59.99">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="" nation="" />
     <RELAY name="vacant" nation="">
      <CLUB name="vacant" nation="" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="" nameprefix="" lastname="" gender="" nation="" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
  <RECORDLIST course="LCM" gender="X" type="WMR" name="Wereld Masters Record" updated="2023-10-31">
   <AGEGROUP agemin="360" agemax="399" calculate="TOTAL" />
   <RECORDS>
    <RECORD swimtime="00:03:36.78">
     <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2013-08-09" nation="" />
     <RELAY name="MISSION VIEJO MASTE" nation="USA">
      <CLUB name="MISSION VIEJO MASTE" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Frank" nameprefix="" lastname="Piemme" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jurgen" nameprefix="" lastname="Schmidt" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:04:19.30">
     <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2013-08-10" nation="" />
     <RELAY name="MISSION VIEJO MASTE" nation="USA">
      <CLUB name="MISSION VIEJO MASTE" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Frank" nameprefix="" lastname="Piemme" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Jurgen" nameprefix="" lastname="Schmidt" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:08:26.02">
     <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2013-07-07" nation="" />
     <RELAY name="MISSION VIEJO NADAD" nation="USA">
      <CLUB name="MISSION VIEJO NADAD" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Frank" nameprefix="" lastname="Piemme" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jurgen" nameprefix="" lastname="Schmidt" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:10:20.46">
     <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
     <MEETINFO city="" date="2013-07-07" nation="" />
     <RELAY name="MISSION VIEJO NADAD" nation="USA">
      <CLUB name="MISSION VIEJO NADAD" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Jurgen" nameprefix="" lastname="Schmidt" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Frank" nameprefix="" lastname="Piemme" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
    <RECORD swimtime="00:18:14.23">
     <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
     <MEETINFO city="" date="2013-07-07" nation="" />
     <RELAY name="MISSION VIEJO NADAD" nation="USA">
      <CLUB name="MISSION VIEJO NADAD" nation="USA" />
      <RELAYPOSITIONS>
       <RELAYPOSITION number="1">
        <ATHLETE firstname="Frank" nameprefix="" lastname="Piemme" gender="M" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="2">
        <ATHLETE firstname="Maurine" nameprefix="" lastname="Kornfeld" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="3">
        <ATHLETE firstname="Rita" nameprefix="" lastname="Simonton" gender="F" nation="USA" />
       </RELAYPOSITION>
       <RELAYPOSITION number="4">
        <ATHLETE firstname="Jurgen" nameprefix="" lastname="Schmidt" gender="M" nation="USA" />
       </RELAYPOSITION>
      </RELAYPOSITIONS>
     </RELAY>
    </RECORD>
   </RECORDS>
  </RECORDLIST>
 </RECORDLISTS>
</LENEX>
